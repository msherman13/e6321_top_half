library verilog;
use verilog.vl_types.all;
entity CLKINVX20TS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end CLKINVX20TS;
