library verilog;
use verilog.vl_types.all;
entity INVXLTS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end INVXLTS;
