##
## LEF for PtnCells ;
## created by First Encounter v08.10-s273_1 on Tue May 14 04:24:54 2013
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MACRO top_level
  CLASS BLOCK ;
  SIZE 5020.0000 BY 2020.0000 ;
  FOREIGN top_level 0 0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 4.32 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.576 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7016 LAYER M3  ;
    ANTENNAMAXAREACAR 2.89563 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 11.3162 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0470146 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2473.7000 0.0000 2473.9000 0.6000 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 50.4189 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 185.523 LAYER MQ  ;
    ANTENNAMAXCUTCAR 4.95496 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2389.2000 0.0000 2389.6000 1.2000 ;
    END
  END reset
  PIN acc_fft_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.66 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.042 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 40.7342 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 156.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2358.1000 0.0000 2358.3000 0.6000 ;
    END
  END acc_fft_get
  PIN acc_fft_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 65.2838 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 248.856 LAYER MQ  ;
    ANTENNAMAXCUTCAR 3.15315 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2429.2000 0.0000 2429.6000 1.2000 ;
    END
  END acc_fft_put
  PIN acc_fir_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.54 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 28.5721 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 113.023 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2325.7000 0.0000 2325.9000 0.6000 ;
    END
  END acc_fir_get
  PIN acc_fir_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.86 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.682 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 9.84 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.296 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 114.608 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 436.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2384.1000 0.0000 2384.3000 0.6000 ;
    END
  END acc_fir_put
  PIN acc_fft_data_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2510.1000 2019.4000 2510.3000 2020.0000 ;
    END
  END acc_fft_data_out[31]
  PIN acc_fft_data_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2510.0000 2018.8000 2510.4000 2020.0000 ;
    END
  END acc_fft_data_out[30]
  PIN acc_fft_data_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2510.9000 2019.4000 2511.1000 2020.0000 ;
    END
  END acc_fft_data_out[29]
  PIN acc_fft_data_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2511.7000 2019.4000 2511.9000 2020.0000 ;
    END
  END acc_fft_data_out[28]
  PIN acc_fft_data_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2511.6000 2018.8000 2512.0000 2020.0000 ;
    END
  END acc_fft_data_out[27]
  PIN acc_fft_data_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2509.3000 2019.4000 2509.5000 2020.0000 ;
    END
  END acc_fft_data_out[26]
  PIN acc_fft_data_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2508.5000 2019.4000 2508.7000 2020.0000 ;
    END
  END acc_fft_data_out[25]
  PIN acc_fft_data_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2508.4000 2018.8000 2508.8000 2020.0000 ;
    END
  END acc_fft_data_out[24]
  PIN acc_fft_data_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2513.3000 2019.4000 2513.5000 2020.0000 ;
    END
  END acc_fft_data_out[23]
  PIN acc_fft_data_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2513.2000 2018.8000 2513.6000 2020.0000 ;
    END
  END acc_fft_data_out[22]
  PIN acc_fft_data_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2506.9000 2019.4000 2507.1000 2020.0000 ;
    END
  END acc_fft_data_out[21]
  PIN acc_fft_data_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2506.8000 2018.8000 2507.2000 2020.0000 ;
    END
  END acc_fft_data_out[20]
  PIN acc_fft_data_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2512.5000 2019.4000 2512.7000 2020.0000 ;
    END
  END acc_fft_data_out[19]
  PIN acc_fft_data_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2514.9000 2019.4000 2515.1000 2020.0000 ;
    END
  END acc_fft_data_out[18]
  PIN acc_fft_data_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2514.8000 2018.8000 2515.2000 2020.0000 ;
    END
  END acc_fft_data_out[17]
  PIN acc_fft_data_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2507.7000 2019.4000 2507.9000 2020.0000 ;
    END
  END acc_fft_data_out[16]
  PIN acc_fft_data_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2505.3000 2019.4000 2505.5000 2020.0000 ;
    END
  END acc_fft_data_out[15]
  PIN acc_fft_data_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2505.2000 2018.8000 2505.6000 2020.0000 ;
    END
  END acc_fft_data_out[14]
  PIN acc_fft_data_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1010.1000 0.6000 1010.3000 ;
    END
  END acc_fft_data_out[13]
  PIN acc_fft_data_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MG ;
        RECT 0.0000 1010.0000 1.2000 1010.4000 ;
    END
  END acc_fft_data_out[12]
  PIN acc_fft_data_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1010.9000 0.6000 1011.1000 ;
    END
  END acc_fft_data_out[11]
  PIN acc_fft_data_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1011.7000 0.6000 1011.9000 ;
    END
  END acc_fft_data_out[10]
  PIN acc_fft_data_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MG ;
        RECT 0.0000 1011.6000 1.2000 1012.0000 ;
    END
  END acc_fft_data_out[9]
  PIN acc_fft_data_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1009.3000 0.6000 1009.5000 ;
    END
  END acc_fft_data_out[8]
  PIN acc_fft_data_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1008.5000 0.6000 1008.7000 ;
    END
  END acc_fft_data_out[7]
  PIN acc_fft_data_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MG ;
        RECT 0.0000 1008.4000 1.2000 1008.8000 ;
    END
  END acc_fft_data_out[6]
  PIN acc_fft_data_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1013.3000 0.6000 1013.5000 ;
    END
  END acc_fft_data_out[5]
  PIN acc_fft_data_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MG ;
        RECT 0.0000 1013.2000 1.2000 1013.6000 ;
    END
  END acc_fft_data_out[4]
  PIN acc_fft_data_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1006.9000 0.6000 1007.1000 ;
    END
  END acc_fft_data_out[3]
  PIN acc_fft_data_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MG ;
        RECT 0.0000 1006.8000 1.2000 1007.2000 ;
    END
  END acc_fft_data_out[2]
  PIN acc_fft_data_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1012.5000 0.6000 1012.7000 ;
    END
  END acc_fft_data_out[1]
  PIN acc_fft_data_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1014.9000 0.6000 1015.1000 ;
    END
  END acc_fft_data_out[0]
  PIN acc_fft_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 36.0045 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2657.7000 0.0000 2657.9000 0.6000 ;
    END
  END acc_fft_data_in[31]
  PIN acc_fft_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.22 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 37.8063 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 140.523 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2662.9000 0.0000 2663.1000 0.6000 ;
    END
  END acc_fft_data_in[30]
  PIN acc_fft_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 21.1396 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 75.5225 LAYER MQ  ;
    ANTENNAMAXCUTCAR 4.95496 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2662.8000 0.0000 2663.2000 1.2000 ;
    END
  END acc_fft_data_in[29]
  PIN acc_fft_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.62 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 42.3108 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 157.189 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2668.5000 0.0000 2668.7000 0.6000 ;
    END
  END acc_fft_data_in[28]
  PIN acc_fft_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.22 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 37.8063 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 140.523 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2604.1000 0.0000 2604.3000 0.6000 ;
    END
  END acc_fft_data_in[27]
  PIN acc_fft_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2613.7000 0.0000 2613.9000 0.6000 ;
    END
  END acc_fft_data_in[26]
  PIN acc_fft_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.02 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 159.914 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 22.7162 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2521.3000 0.0000 2521.5000 0.6000 ;
    END
  END acc_fft_data_in[25]
  PIN acc_fft_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.978 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 29.0225 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 116.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2526.1000 0.0000 2526.3000 0.6000 ;
    END
  END acc_fft_data_in[24]
  PIN acc_fft_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.34 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 27.8964 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 103.856 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2604.9000 0.0000 2605.1000 0.6000 ;
    END
  END acc_fft_data_in[23]
  PIN acc_fft_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.62 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 42.3108 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 157.189 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2675.3000 0.0000 2675.5000 0.6000 ;
    END
  END acc_fft_data_in[22]
  PIN acc_fft_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2666.5000 0.0000 2666.7000 0.6000 ;
    END
  END acc_fft_data_in[21]
  PIN acc_fft_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2608.9000 0.0000 2609.1000 0.6000 ;
    END
  END acc_fft_data_in[20]
  PIN acc_fft_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 54.9234 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 208.856 LAYER MQ  ;
    ANTENNAMAXCUTCAR 3.15315 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2521.2000 0.0000 2521.6000 1.2000 ;
    END
  END acc_fft_data_in[19]
  PIN acc_fft_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.62 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 42.3108 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 157.189 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2572.5000 0.0000 2572.7000 0.6000 ;
    END
  END acc_fft_data_in[18]
  PIN acc_fft_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.25 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 39.3829 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 149.689 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2535.7000 0.0000 2535.9000 0.6000 ;
    END
  END acc_fft_data_in[17]
  PIN acc_fft_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 119.563 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 446.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2546.9000 0.0000 2547.1000 0.6000 ;
    END
  END acc_fft_data_in[16]
  PIN acc_fft_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.38 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 39.6081 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 147.189 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2598.9000 0.0000 2599.1000 0.6000 ;
    END
  END acc_fft_data_in[15]
  PIN acc_fft_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2570.9000 0.0000 2571.1000 0.6000 ;
    END
  END acc_fft_data_in[14]
  PIN acc_fft_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2621.3000 0.0000 2621.5000 0.6000 ;
    END
  END acc_fft_data_in[13]
  PIN acc_fft_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2566.1000 0.0000 2566.3000 0.6000 ;
    END
  END acc_fft_data_in[12]
  PIN acc_fft_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 58.527 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 217.189 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2670.9000 0.0000 2671.1000 0.6000 ;
    END
  END acc_fft_data_in[11]
  PIN acc_fft_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 36.0045 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2673.7000 0.0000 2673.9000 0.6000 ;
    END
  END acc_fft_data_in[10]
  PIN acc_fft_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.34 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 27.8964 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 103.856 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2663.7000 0.0000 2663.9000 0.6000 ;
    END
  END acc_fft_data_in[9]
  PIN acc_fft_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.78 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.834 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 55.3739 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 207.189 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2658.5000 0.0000 2658.7000 0.6000 ;
    END
  END acc_fft_data_in[8]
  PIN acc_fft_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 74.2928 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 285.523 LAYER MQ  ;
    ANTENNAMAXCUTCAR 3.15315 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2535.6000 0.0000 2536.0000 1.2000 ;
    END
  END acc_fft_data_in[7]
  PIN acc_fft_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 36.0045 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2566.9000 0.0000 2567.1000 0.6000 ;
    END
  END acc_fft_data_in[6]
  PIN acc_fft_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 31.5 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 112.189 LAYER MQ  ;
    ANTENNAMAXCUTCAR 4.95496 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2598.8000 0.0000 2599.2000 1.2000 ;
    END
  END acc_fft_data_in[5]
  PIN acc_fft_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.22 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.514 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 24.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.648 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2136 LAYER M3  ;
    ANTENNAMAXAREACAR 116.96 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 438.586 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.561798 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2527.7000 0.0000 2527.9000 0.6000 ;
    END
  END acc_fft_data_in[4]
  PIN acc_fft_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2636.1000 0.0000 2636.3000 0.6000 ;
    END
  END acc_fft_data_in[3]
  PIN acc_fft_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.722 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 3.08 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.136 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 39.3829 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 156.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2560.9000 0.0000 2561.1000 0.6000 ;
    END
  END acc_fft_data_in[2]
  PIN acc_fft_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.65 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 52.2207 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 193.856 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2584.1000 0.0000 2584.3000 0.6000 ;
    END
  END acc_fft_data_in[1]
  PIN acc_fft_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.78 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 16.8604 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 66.3559 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2664.5000 0.0000 2664.7000 0.6000 ;
    END
  END acc_fft_data_in[0]
  PIN acc_fir_data_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MG ;
        RECT 0.0000 1014.8000 1.2000 1015.2000 ;
    END
  END acc_fir_data_out[31]
  PIN acc_fir_data_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1007.7000 0.6000 1007.9000 ;
    END
  END acc_fir_data_out[30]
  PIN acc_fir_data_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1005.3000 0.6000 1005.5000 ;
    END
  END acc_fir_data_out[29]
  PIN acc_fir_data_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MG ;
        RECT 0.0000 1005.2000 1.2000 1005.6000 ;
    END
  END acc_fir_data_out[28]
  PIN acc_fir_data_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2516.5000 2019.4000 2516.7000 2020.0000 ;
    END
  END acc_fir_data_out[27]
  PIN acc_fir_data_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2503.6000 2018.8000 2504.0000 2020.0000 ;
    END
  END acc_fir_data_out[26]
  PIN acc_fir_data_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2514.1000 2019.4000 2514.3000 2020.0000 ;
    END
  END acc_fir_data_out[25]
  PIN acc_fir_data_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2518.0000 2018.8000 2518.4000 2020.0000 ;
    END
  END acc_fir_data_out[24]
  PIN acc_fir_data_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2506.1000 2019.4000 2506.3000 2020.0000 ;
    END
  END acc_fir_data_out[23]
  PIN acc_fir_data_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2502.0000 2018.8000 2502.4000 2020.0000 ;
    END
  END acc_fir_data_out[22]
  PIN acc_fir_data_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2519.6000 2018.8000 2520.0000 2020.0000 ;
    END
  END acc_fir_data_out[21]
  PIN acc_fir_data_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2500.4000 2018.8000 2500.8000 2020.0000 ;
    END
  END acc_fir_data_out[20]
  PIN acc_fir_data_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2515.7000 2019.4000 2515.9000 2020.0000 ;
    END
  END acc_fir_data_out[19]
  PIN acc_fir_data_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2521.2000 2018.8000 2521.6000 2020.0000 ;
    END
  END acc_fir_data_out[18]
  PIN acc_fir_data_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2504.5000 2019.4000 2504.7000 2020.0000 ;
    END
  END acc_fir_data_out[17]
  PIN acc_fir_data_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2498.8000 2018.8000 2499.2000 2020.0000 ;
    END
  END acc_fir_data_out[16]
  PIN acc_fir_data_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2516.4000 2018.8000 2516.8000 2020.0000 ;
    END
  END acc_fir_data_out[15]
  PIN acc_fir_data_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2522.8000 2018.8000 2523.2000 2020.0000 ;
    END
  END acc_fir_data_out[14]
  PIN acc_fir_data_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2503.7000 2019.4000 2503.9000 2020.0000 ;
    END
  END acc_fir_data_out[13]
  PIN acc_fir_data_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2497.2000 2018.8000 2497.6000 2020.0000 ;
    END
  END acc_fir_data_out[12]
  PIN acc_fir_data_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2517.3000 2019.4000 2517.5000 2020.0000 ;
    END
  END acc_fir_data_out[11]
  PIN acc_fir_data_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2524.4000 2018.8000 2524.8000 2020.0000 ;
    END
  END acc_fir_data_out[10]
  PIN acc_fir_data_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2502.9000 2019.4000 2503.1000 2020.0000 ;
    END
  END acc_fir_data_out[9]
  PIN acc_fir_data_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2495.6000 2018.8000 2496.0000 2020.0000 ;
    END
  END acc_fir_data_out[8]
  PIN acc_fir_data_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2518.1000 2019.4000 2518.3000 2020.0000 ;
    END
  END acc_fir_data_out[7]
  PIN acc_fir_data_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2526.0000 2018.8000 2526.4000 2020.0000 ;
    END
  END acc_fir_data_out[6]
  PIN acc_fir_data_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2502.1000 2019.4000 2502.3000 2020.0000 ;
    END
  END acc_fir_data_out[5]
  PIN acc_fir_data_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2494.0000 2018.8000 2494.4000 2020.0000 ;
    END
  END acc_fir_data_out[4]
  PIN acc_fir_data_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2518.9000 2019.4000 2519.1000 2020.0000 ;
    END
  END acc_fir_data_out[3]
  PIN acc_fir_data_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2527.6000 2018.8000 2528.0000 2020.0000 ;
    END
  END acc_fir_data_out[2]
  PIN acc_fir_data_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2501.3000 2019.4000 2501.5000 2020.0000 ;
    END
  END acc_fir_data_out[1]
  PIN acc_fir_data_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 2492.4000 2018.8000 2492.8000 2020.0000 ;
    END
  END acc_fir_data_out[0]
  PIN acc_fir_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 100.714 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 16.8604 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 66.3559 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2296.5000 0.0000 2296.7000 0.6000 ;
    END
  END acc_fir_data_in[31]
  PIN acc_fir_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.26 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 8.88 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.448 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 108.302 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 409.689 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2286.1000 0.0000 2286.3000 0.6000 ;
    END
  END acc_fir_data_in[30]
  PIN acc_fir_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.586 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 4.88 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.352 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 65.0586 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 246.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2301.3000 0.0000 2301.5000 0.6000 ;
    END
  END acc_fir_data_in[29]
  PIN acc_fir_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.98 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.826 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 6.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.456 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 98.8423 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 373.023 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2305.7000 0.0000 2305.9000 0.6000 ;
    END
  END acc_fir_data_in[28]
  PIN acc_fir_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 155.824 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 582.189 LAYER MQ  ;
    ANTENNAMAXCUTCAR 2.7027 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2296.4000 0.0000 2296.8000 1.2000 ;
    END
  END acc_fir_data_in[27]
  PIN acc_fir_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 47.7162 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 175.523 LAYER MQ  ;
    ANTENNAMAXCUTCAR 4.95496 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2301.2000 0.0000 2301.6000 1.2000 ;
    END
  END acc_fir_data_in[26]
  PIN acc_fir_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.018 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 9 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.04 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 107.851 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 409.689 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2295.7000 0.0000 2295.9000 0.6000 ;
    END
  END acc_fir_data_in[25]
  PIN acc_fir_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 42.0856 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 163.023 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2298.1000 0.0000 2298.3000 0.6000 ;
    END
  END acc_fir_data_in[24]
  PIN acc_fir_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.62 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 42.3108 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 157.189 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2586.5000 0.0000 2586.7000 0.6000 ;
    END
  END acc_fir_data_in[23]
  PIN acc_fir_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 58.527 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 217.189 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2677.3000 0.0000 2677.5000 0.6000 ;
    END
  END acc_fir_data_in[22]
  PIN acc_fir_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.22 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.314 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 60.3288 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 223.856 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2599.7000 0.0000 2599.9000 0.6000 ;
    END
  END acc_fir_data_in[21]
  PIN acc_fir_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 36.0045 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2580.9000 0.0000 2581.1000 0.6000 ;
    END
  END acc_fir_data_in[20]
  PIN acc_fir_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.778 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 4.24775 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 19.6892 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2545.3000 0.0000 2545.5000 0.6000 ;
    END
  END acc_fir_data_in[19]
  PIN acc_fir_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.22 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 37.8063 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 140.523 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2609.7000 0.0000 2609.9000 0.6000 ;
    END
  END acc_fir_data_in[18]
  PIN acc_fir_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2582.5000 0.0000 2582.7000 0.6000 ;
    END
  END acc_fir_data_in[17]
  PIN acc_fir_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2593.3000 0.0000 2593.5000 0.6000 ;
    END
  END acc_fir_data_in[16]
  PIN acc_fir_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 42.3108 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 152.189 LAYER MQ  ;
    ANTENNAMAXCUTCAR 4.95496 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2677.2000 0.0000 2677.6000 1.2000 ;
    END
  END acc_fir_data_in[15]
  PIN acc_fir_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.66 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.642 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 76.545 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 283.856 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2691.7000 0.0000 2691.9000 0.6000 ;
    END
  END acc_fir_data_in[14]
  PIN acc_fir_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2623.7000 0.0000 2623.9000 0.6000 ;
    END
  END acc_fir_data_in[13]
  PIN acc_fir_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 58.527 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 217.189 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2692.5000 0.0000 2692.7000 0.6000 ;
    END
  END acc_fir_data_in[12]
  PIN acc_fir_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.0946 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2647.3000 0.0000 2647.5000 0.6000 ;
    END
  END acc_fir_data_in[11]
  PIN acc_fir_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.26 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2  ;
    ANTENNAMAXAREACAR 26.9955 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 100.523 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2676.1000 0.0000 2676.3000 0.6000 ;
    END
  END acc_fir_data_in[10]
  PIN acc_fir_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ  ;
    ANTENNAMAXAREACAR 31.5 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 112.189 LAYER MQ  ;
    ANTENNAMAXCUTCAR 4.95496 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2658.0000 0.0000 2658.4000 1.2000 ;
    END
  END acc_fir_data_in[9]
  PIN acc_fir_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 14.1577 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 56.3559 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2659.7000 0.0000 2659.9000 0.6000 ;
    END
  END acc_fir_data_in[8]
  PIN acc_fir_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 111.005 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 416.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2417.3000 0.0000 2417.5000 0.6000 ;
    END
  END acc_fir_data_in[7]
  PIN acc_fir_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 6.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.456 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 96.5901 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 366.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2379.3000 0.0000 2379.5000 0.6000 ;
    END
  END acc_fir_data_in[6]
  PIN acc_fir_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 3.4 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.32 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 41.1847 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 163.023 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2380.1000 0.0000 2380.3000 0.6000 ;
    END
  END acc_fir_data_in[5]
  PIN acc_fir_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.86 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.882 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1056 LAYER M3  ;
    ANTENNAMAXAREACAR 61.5417 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 231.644 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.51515 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2435.7000 0.0000 2435.9000 0.6000 ;
    END
  END acc_fir_data_in[4]
  PIN acc_fir_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.58 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.546 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 143.887 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 536.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2482.5000 0.0000 2482.7000 0.6000 ;
    END
  END acc_fir_data_in[3]
  PIN acc_fir_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.33 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 3.44 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.32 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 56.9505 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 219.689 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2448.5000 0.0000 2448.7000 0.6000 ;
    END
  END acc_fir_data_in[2]
  PIN acc_fir_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.578 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 47.0405 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 179.689 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2498.5000 0.0000 2498.7000 0.6000 ;
    END
  END acc_fir_data_in[1]
  PIN acc_fir_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.74 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.938 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 70.464 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 266.356 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2496.5000 0.0000 2496.7000 0.6000 ;
    END
  END acc_fir_data_in[0]
  PIN fft_enable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7272 LAYER MQ  ;
    ANTENNAMAXAREACAR 23.6574 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 88.4455 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.892307 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2418.8000 0.0000 2419.2000 1.2000 ;
    END
  END fft_enable
  PIN fir_enable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.34 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.706 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M2  ;
    ANTENNAMAXAREACAR 133.833 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 496.976 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2  ;
    ANTENNAMAXCUTCAR 1.6129 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 13.28 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.728 LAYER M3  ;
    ANTENNAGATEAREA 4.1152 LAYER M3  ;
    ANTENNAMAXAREACAR 137.06 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 509.06 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2322.1000 0.0000 2322.3000 0.6000 ;
    END
  END fir_enable
  PIN to_fft_empty
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 16.44 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.16 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.5808 LAYER M3  ;
    ANTENNAMAXAREACAR 13.8147 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 52.3224 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.806452 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2356.9000 0.0000 2357.1000 0.6000 ;
    END
  END to_fft_empty
  PIN from_fft_full
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.62 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.994 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M3  ;
    ANTENNAMAXAREACAR 2.62364 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 9.56523 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2414.5000 0.0000 2414.7000 0.6000 ;
    END
  END from_fft_full
  PIN to_fir_empty
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.01 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 8.04 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.5328 LAYER M3  ;
    ANTENNAMAXAREACAR 92.242 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 340.974 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.98413 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2316.1000 0.0000 2316.3000 0.6000 ;
    END
  END to_fir_empty
  PIN from_fir_full
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER MQ  ;
    ANTENNAMAXAREACAR 4.68432 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 17.0706 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.136364 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2383.6000 0.0000 2384.0000 1.2000 ;
    END
  END from_fir_full
  PIN ram_read_enable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.207 LAYER MQ  ;
    ANTENNAMAXAREACAR 1.55162 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 5.29591 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.0666019 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2325.2000 0.0000 2325.6000 1.2000 ;
    END
  END ram_read_enable
  PIN ram_write_enable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.898 LAYER M2  ;
    ANTENNAMAXAREACAR 0.938854 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 3.46253 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0138026 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2331.3000 0.0000 2331.5000 0.6000 ;
    END
  END ram_write_enable
  PIN addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.66 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.642 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 20.04 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.184 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 2.90451 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 10.7408 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2394.1000 0.0000 2394.3000 0.6000 ;
    END
  END addr[31]
  PIN addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.38 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.106 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 14.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.76 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.38214 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.02438 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2389.3000 0.0000 2389.5000 0.6000 ;
    END
  END addr[30]
  PIN addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.178 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 17.32 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.824 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.98029 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 7.24375 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2392.1000 0.0000 2392.3000 0.6000 ;
    END
  END addr[29]
  PIN addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.38 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.906 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 14.8 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.056 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.52311 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.48796 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2399.7000 0.0000 2399.9000 0.6000 ;
    END
  END addr[28]
  PIN addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.02 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.474 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 3.69711 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 13.4747 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 12.28 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.88 LAYER M3  ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 4.28931 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 15.6872 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0617284 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2405.7000 0.0000 2405.9000 0.6000 ;
    END
  END addr[27]
  PIN addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER MQ  ;
    ANTENNAMAXAREACAR 3.96813 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 14.5488 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.108025 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2399.6000 0.0000 2400.0000 1.2000 ;
    END
  END addr[26]
  PIN addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 12.84 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.248 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 4.40312 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 16.2083 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2403.7000 0.0000 2403.9000 0.6000 ;
    END
  END addr[25]
  PIN addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 17.4 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.416 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.64988 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 6.06605 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2404.5000 0.0000 2404.7000 0.6000 ;
    END
  END addr[24]
  PIN addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER MQ  ;
    ANTENNAMAXAREACAR 1.29244 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 4.77197 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.100309 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2417.2000 0.0000 2417.6000 1.2000 ;
    END
  END addr[23]
  PIN addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.922 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 15.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.72 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.42303 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.14514 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2415.7000 0.0000 2415.9000 0.6000 ;
    END
  END addr[22]
  PIN addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.74 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 10.52 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.072 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.14309 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 4.07477 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0578704 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2429.3000 0.0000 2429.5000 0.6000 ;
    END
  END addr[21]
  PIN addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.866 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.97257 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 7.22234 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 8.44 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER M3  ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 2.37959 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 8.74973 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2436.9000 0.0000 2437.1000 0.6000 ;
    END
  END addr[20]
  PIN addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.38 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.106 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 16.04 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.088 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.82967 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 6.68642 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2439.7000 0.0000 2439.9000 0.6000 ;
    END
  END addr[19]
  PIN addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 15.48 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.016 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 2.19248 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 8.02886 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2427.3000 0.0000 2427.5000 0.6000 ;
    END
  END addr[18]
  PIN addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.466 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 18 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.192 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 2.00058 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 7.32994 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2434.1000 0.0000 2434.3000 0.6000 ;
    END
  END addr[17]
  PIN addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.42 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.65 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.912 LAYER M2  ;
    ANTENNAMAXAREACAR 0.858565 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 3.01487 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2  ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 18.44 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.672 LAYER M3  ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.74784 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 6.3266 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2428.5000 0.0000 2428.7000 0.6000 ;
    END
  END addr[16]
  PIN addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.22 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.514 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 17.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.712 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 2.05035 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 7.5294 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2432.9000 0.0000 2433.1000 0.6000 ;
    END
  END addr[15]
  PIN addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER MQ  ;
    ANTENNAMAXAREACAR 2.26408 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 8.29271 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.100309 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2435.6000 0.0000 2436.0000 1.2000 ;
    END
  END addr[14]
  PIN addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.66 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 12.48 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.768 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.60613 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.87253 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2437.7000 0.0000 2437.9000 0.6000 ;
    END
  END addr[13]
  PIN addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.42 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.202 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.78738 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 6.4515 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 14.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.352 LAYER M3  ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 2.49919 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 9.12087 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2434.9000 0.0000 2435.1000 0.6000 ;
    END
  END addr[12]
  PIN addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER MQ  ;
    ANTENNAMAXAREACAR 3.00887 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 11.0586 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.123457 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2427.6000 0.0000 2428.0000 1.2000 ;
    END
  END addr[11]
  PIN addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 13.24 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.432 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.27334 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 4.72577 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2420.5000 0.0000 2420.7000 0.6000 ;
    END
  END addr[10]
  PIN addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.29 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 15.84 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.2 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 3.11262 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 11.4262 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2418.1000 0.0000 2418.3000 0.6000 ;
    END
  END addr[9]
  PIN addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.62 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.994 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 17.56 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.416 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 3.61223 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 13.2677 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2419.3000 0.0000 2419.5000 0.6000 ;
    END
  END addr[8]
  PIN addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.58 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 18.24 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.376 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 2.28669 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 8.39259 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2413.7000 0.0000 2413.9000 0.6000 ;
    END
  END addr[7]
  PIN addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 19.56 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.112 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.8684 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 6.78696 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2412.1000 0.0000 2412.3000 0.6000 ;
    END
  END addr[6]
  PIN addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.56 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.12 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 17.56 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.008 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.91107 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 7.00085 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2402.9000 0.0000 2403.1000 0.6000 ;
    END
  END addr[5]
  PIN addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.33 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 18.4 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.968 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 3.3532 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 12.5568 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2411.3000 0.0000 2411.5000 0.6000 ;
    END
  END addr[4]
  PIN addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.42 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.554 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 19.4 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.224 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.64834 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.95841 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2398.5000 0.0000 2398.7000 0.6000 ;
    END
  END addr[3]
  PIN addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.34 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.106 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 17.28 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.232 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.28067 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 4.63164 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0578704 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2400.9000 0.0000 2401.1000 0.6000 ;
    END
  END addr[2]
  PIN addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.74 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.338 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 13.08 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.136 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.81424 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 6.5865 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2401.7000 0.0000 2401.9000 0.6000 ;
    END
  END addr[1]
  PIN addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 16.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.456 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3  ;
    ANTENNAMAXAREACAR 1.85783 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 6.75085 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2406.5000 0.0000 2406.7000 0.6000 ;
    END
  END addr[0]
  PIN data_bus[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.38 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.6 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 2.49363 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 9.1706 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2514.9000 0.0000 2515.1000 0.6000 ;
    END
  END data_bus[31]
  PIN data_bus[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.42 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.354 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 3.88 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.948 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 2.29688 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 8.52824 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2515.7000 0.0000 2515.9000 0.6000 ;
    END
  END data_bus[30]
  PIN data_bus[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.978 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 1.82002 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 6.70069 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2524.5000 0.0000 2524.7000 0.6000 ;
    END
  END data_bus[29]
  PIN data_bus[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.02 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.074 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 1.20289 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 4.37454 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2520.1000 0.0000 2520.3000 0.6000 ;
    END
  END data_bus[28]
  PIN data_bus[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.66 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.738 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 6.3397 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 23.3888 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2505.7000 0.0000 2505.9000 0.6000 ;
    END
  END data_bus[27]
  PIN data_bus[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.418 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 5.17859 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 18.9561 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2532.1000 0.0000 2532.3000 0.6000 ;
    END
  END data_bus[26]
  PIN data_bus[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.02 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.474 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 3.93762 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 14.469 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2508.5000 0.0000 2508.7000 0.6000 ;
    END
  END data_bus[25]
  PIN data_bus[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.02 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.474 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.6 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 1.69271 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 6.23773 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2490.9000 0.0000 2491.1000 0.6000 ;
    END
  END data_bus[24]
  PIN data_bus[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.26 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.762 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.45174 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 5.16678 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2597.7000 0.0000 2597.9000 0.6000 ;
    END
  END data_bus[23]
  PIN data_bus[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.66 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.4022 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 5.06701 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2624.9000 0.0000 2625.1000 0.6000 ;
    END
  END data_bus[22]
  PIN data_bus[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.54 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.2434 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 4.39595 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2607.7000 0.0000 2607.9000 0.6000 ;
    END
  END data_bus[21]
  PIN data_bus[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.98 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.426 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.66007 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 5.93762 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2602.5000 0.0000 2602.7000 0.6000 ;
    END
  END data_bus[20]
  PIN data_bus[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 4.89641 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 18.0711 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2547.7000 0.0000 2547.9000 0.6000 ;
    END
  END data_bus[19]
  PIN data_bus[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.09 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.8684 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 6.70845 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2569.3000 0.0000 2569.5000 0.6000 ;
    END
  END data_bus[18]
  PIN data_bus[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.38 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 3.92 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 2.37326 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 8.73542 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2538.1000 0.0000 2538.3000 0.6000 ;
    END
  END data_bus[17]
  PIN data_bus[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.82 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.834 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.12 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 2.63808 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 9.68472 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2533.7000 0.0000 2533.9000 0.6000 ;
    END
  END data_bus[16]
  PIN data_bus[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.82 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.434 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.03507 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 3.62512 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2612.1000 0.0000 2612.3000 0.6000 ;
    END
  END data_bus[15]
  PIN data_bus[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.26 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.762 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.45174 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 5.16678 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2588.9000 0.0000 2589.1000 0.6000 ;
    END
  END data_bus[14]
  PIN data_bus[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 0.826736 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 2.85428 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2616.9000 0.0000 2617.1000 0.6000 ;
    END
  END data_bus[13]
  PIN data_bus[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ  ;
    ANTENNAMAXAREACAR 0.629977 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 2.04063 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2582.0000 0.0000 2582.4000 1.2000 ;
    END
  END data_bus[12]
  PIN data_bus[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 0.826736 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 2.85428 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2626.1000 0.0000 2626.3000 0.6000 ;
    END
  END data_bus[11]
  PIN data_bus[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.34 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.058 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 1.52488 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 5.43738 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2619.7000 0.0000 2619.9000 0.6000 ;
    END
  END data_bus[10]
  PIN data_bus[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2  ;
    ANTENNAMAXAREACAR 0.826736 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 2.85428 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 2634.1000 0.0000 2634.3000 0.6000 ;
    END
  END data_bus[9]
  PIN data_bus[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ  ;
    ANTENNAMAXAREACAR 1.19711 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 4.09618 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2625.2000 0.0000 2625.6000 1.2000 ;
    END
  END data_bus[8]
  PIN data_bus[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.73 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 4.07234 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 15.0016 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2500.5000 0.0000 2500.7000 0.6000 ;
    END
  END data_bus[7]
  PIN data_bus[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ  ;
    ANTENNAMAXAREACAR 1.00174 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 3.66076 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2514.8000 0.0000 2515.2000 1.2000 ;
    END
  END data_bus[6]
  PIN data_bus[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ  ;
    ANTENNAMAXAREACAR 2.23877 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 8.20729 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2496.4000 0.0000 2496.8000 1.2000 ;
    END
  END data_bus[5]
  PIN data_bus[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.74 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 4 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.392 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 1.43438 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.31667 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2516.5000 0.0000 2516.7000 0.6000 ;
    END
  END data_bus[4]
  PIN data_bus[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.52 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 2.17419 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 7.97847 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2539.3000 0.0000 2539.5000 0.6000 ;
    END
  END data_bus[3]
  PIN data_bus[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ  ;
    ANTENNAMAXAREACAR 3.211 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 11.6332 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2516.4000 0.0000 2516.8000 1.2000 ;
    END
  END data_bus[2]
  PIN data_bus[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ  ;
    ANTENNAMAXAREACAR 6.19711 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 22.5962 LAYER MQ  ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VQ  ;
    PORT
      LAYER MQ ;
        RECT 2508.4000 0.0000 2508.8000 1.2000 ;
    END
  END data_bus[1]
  PIN data_bus[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3  ;
    ANTENNAMAXAREACAR 4.03854 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 14.8236 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 2530.1000 0.0000 2530.3000 0.6000 ;
    END
  END data_bus[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power strip data as pin
    PORT
    END
# end of P/G power strip data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power strip data as pin
    PORT
    END
# end of P/G power strip data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 5020.0000 2020.0000 ;
    LAYER M2 ;
      RECT 2521.0200 2017.4800 5020.0000 2020.0000 ;
      RECT 0.0000 2017.4800 2499.3800 2020.0000 ;
      RECT 0.0000 2.5200 5020.0000 2017.4800 ;
      RECT 2694.6200 0.0000 5020.0000 2.5200 ;
      RECT 2679.4200 0.0000 2689.7800 2.5200 ;
      RECT 2649.4200 0.0000 2655.7800 2.5200 ;
      RECT 2638.2200 0.0000 2645.3800 2.5200 ;
      RECT 2628.2200 0.0000 2632.1800 2.5200 ;
      RECT 2595.4200 0.0000 2595.7800 2.5200 ;
      RECT 2591.0200 0.0000 2591.3800 2.5200 ;
      RECT 2574.6200 0.0000 2578.9800 2.5200 ;
      RECT 2563.0200 0.0000 2564.1800 2.5200 ;
      RECT 2549.8200 0.0000 2558.9800 2.5200 ;
      RECT 2541.4200 0.0000 2543.3800 2.5200 ;
      RECT 2510.6200 0.0000 2512.9800 2.5200 ;
      RECT 2502.6200 0.0000 2503.7800 2.5200 ;
      RECT 2493.0200 0.0000 2494.5800 2.5200 ;
      RECT 2484.6200 0.0000 2488.9800 2.5200 ;
      RECT 2475.8200 0.0000 2480.5800 2.5200 ;
      RECT 2450.6200 0.0000 2471.7800 2.5200 ;
      RECT 2441.8200 0.0000 2446.5800 2.5200 ;
      RECT 2422.6200 0.0000 2425.3800 2.5200 ;
      RECT 2408.6200 0.0000 2409.3800 2.5200 ;
      RECT 2396.2200 0.0000 2396.5800 2.5200 ;
      RECT 2386.2200 0.0000 2387.3800 2.5200 ;
      RECT 2360.2200 0.0000 2377.3800 2.5200 ;
      RECT 2333.4200 0.0000 2354.9800 2.5200 ;
      RECT 2327.8200 0.0000 2329.3800 2.5200 ;
      RECT 2318.2200 0.0000 2320.1800 2.5200 ;
      RECT 2307.8200 0.0000 2314.1800 2.5200 ;
      RECT 2303.4200 0.0000 2303.7800 2.5200 ;
      RECT 2288.2200 0.0000 2293.7800 2.5200 ;
      RECT 0.0000 0.0000 2284.1800 2.5200 ;
    LAYER M3 ;
      RECT 0.0000 1017.0200 5020.0000 2020.0000 ;
      RECT 2.5200 1012.9800 5020.0000 1017.0200 ;
      RECT 2.5200 1011.3800 5020.0000 1012.9800 ;
      RECT 2.5200 1010.5800 5020.0000 1011.3800 ;
      RECT 2.5200 1009.7800 5020.0000 1010.5800 ;
      RECT 2.5200 1008.9800 5020.0000 1009.7800 ;
      RECT 2.5200 1008.1800 5020.0000 1008.9800 ;
      RECT 2.5200 1007.3800 5020.0000 1008.1800 ;
      RECT 2.5200 1006.5800 5020.0000 1007.3800 ;
      RECT 2.5200 1005.7800 5020.0000 1006.5800 ;
      RECT 2.5200 1004.9800 5020.0000 1005.7800 ;
      RECT 2.5200 1003.3800 5020.0000 1004.9800 ;
      RECT 0.0000 0.0000 5020.0000 1003.3800 ;
    LAYER MQ ;
      RECT 2529.9200 2016.8800 5020.0000 2020.0000 ;
      RECT 0.0000 2016.8800 2490.4800 2020.0000 ;
      RECT 0.0000 3.1200 5020.0000 2016.8800 ;
      RECT 2679.5200 0.0000 5020.0000 3.1200 ;
      RECT 2665.1200 0.0000 2675.2800 3.1200 ;
      RECT 2660.3200 0.0000 2660.8800 3.1200 ;
      RECT 2627.5200 0.0000 2656.0800 3.1200 ;
      RECT 2601.1200 0.0000 2623.2800 3.1200 ;
      RECT 2584.3200 0.0000 2596.8800 3.1200 ;
      RECT 2537.9200 0.0000 2580.0800 3.1200 ;
      RECT 2523.5200 0.0000 2533.6800 3.1200 ;
      RECT 2518.7200 0.0000 2519.2800 3.1200 ;
      RECT 2510.7200 0.0000 2512.8800 3.1200 ;
      RECT 2498.7200 0.0000 2506.4800 3.1200 ;
      RECT 2437.9200 0.0000 2494.4800 3.1200 ;
      RECT 2431.5200 0.0000 2433.6800 3.1200 ;
      RECT 2421.1200 0.0000 2425.6800 3.1200 ;
      RECT 2401.9200 0.0000 2415.2800 3.1200 ;
      RECT 2391.5200 0.0000 2397.6800 3.1200 ;
      RECT 2385.9200 0.0000 2387.2800 3.1200 ;
      RECT 2327.5200 0.0000 2381.6800 3.1200 ;
      RECT 2303.5200 0.0000 2323.2800 3.1200 ;
      RECT 2298.7200 0.0000 2299.2800 3.1200 ;
      RECT 0.0000 0.0000 2294.4800 3.1200 ;
  END
END top_level

END LIBRARY
