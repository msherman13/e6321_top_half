library verilog;
use verilog.vl_types.all;
entity DLY3X4TS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end DLY3X4TS;
