library verilog;
use verilog.vl_types.all;
entity INVX12TS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end INVX12TS;
