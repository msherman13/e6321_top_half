library verilog;
use verilog.vl_types.all;
entity HOLDX1TS is
    port(
        Y               : inout  vl_logic
    );
end HOLDX1TS;
