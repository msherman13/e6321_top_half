library verilog;
use verilog.vl_types.all;
entity CLKBUFX12TS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end CLKBUFX12TS;
