library verilog;
use verilog.vl_types.all;
entity top_level_tb is
end top_level_tb;
