library verilog;
use verilog.vl_types.all;
entity udp_sedff is
    // This module cannot be connected to from
    // VHDL because it has unnamed ports.
end udp_sedff;
