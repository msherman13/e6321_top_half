library verilog;
use verilog.vl_types.all;
entity RFRDX1TS is
    port(
        BRB             : out    vl_logic;
        RB              : in     vl_logic
    );
end RFRDX1TS;
