library verilog;
use verilog.vl_types.all;
entity BUFX16TS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end BUFX16TS;
