
module dc_router_top ( chipselect, clk, reset, instruction, offset, filesize, 
        acc_done, fft_enable, fir_enable, iir_enable, data_bus, fft_data_in, 
        fir_data_in, iir_data_in, fft_data_out, fir_data_out, iir_data_out, 
        to_fft_empty, to_fft_full, from_fft_empty, from_fft_full, to_fir_empty, 
        to_fir_full, from_fir_empty, from_fir_full, to_iir_empty, to_iir_full, 
        from_iir_empty, from_iir_full, fft_put_req, fft_get_req, fir_put_req, 
        fir_get_req, iir_put_req, iir_get_req, ram_read_enable, 
        ram_write_enable, addr );
  input [31:0] instruction;
  input [31:0] offset;
  input [31:0] filesize;
  inout [31:0] data_bus;
  input [31:0] fft_data_in;
  input [31:0] fir_data_in;
  input [31:0] iir_data_in;
  output [31:0] fft_data_out;
  output [31:0] fir_data_out;
  output [31:0] iir_data_out;
  output [31:0] addr;
  input chipselect, clk, reset, to_fft_empty, to_fft_full, from_fft_empty,
         from_fft_full, to_fir_empty, to_fir_full, from_fir_empty,
         from_fir_full, to_iir_empty, to_iir_full, from_iir_empty,
         from_iir_full;
  output acc_done, fft_enable, fir_enable, iir_enable, fft_put_req,
         fft_get_req, fir_put_req, fir_get_req, iir_put_req, iir_get_req,
         ram_read_enable, ram_write_enable;
  wire   n2814, n2815, data_to_fft, data_from_fft, data_to_fir, data_from_fir,
         data_to_iir, data_from_iir, fft_read_done, fir_read_done,
         fir_write_done, iir_read_done, iir_write_done, fft_put_req_reg,
         fir_put_req_reg, fir_get_req_reg, iir_put_req_reg, iir_get_req_reg,
         \pla_top/N59 , \pla_top/instruction_valid , \addr_calc/N224 ,
         \addr_calc/N223 , \addr_calc/N220 , \addr_calc/N219 ,
         \addr_calc/N217 , \addr_calc/N216 , \addr_calc/iir_write_addr[31] ,
         \addr_calc/iir_write_addr[30] , \addr_calc/iir_write_addr[29] ,
         \addr_calc/iir_write_addr[28] , \addr_calc/iir_write_addr[27] ,
         \addr_calc/iir_write_addr[26] , \addr_calc/iir_write_addr[25] ,
         \addr_calc/iir_write_addr[24] , \addr_calc/iir_write_addr[23] ,
         \addr_calc/iir_write_addr[22] , \addr_calc/iir_write_addr[21] ,
         \addr_calc/iir_write_addr[20] , \addr_calc/iir_write_addr[19] ,
         \addr_calc/iir_write_addr[18] , \addr_calc/iir_write_addr[17] ,
         \addr_calc/iir_write_addr[16] , \addr_calc/iir_write_addr[15] ,
         \addr_calc/iir_write_addr[14] , \addr_calc/iir_write_addr[13] ,
         \addr_calc/iir_write_addr[12] , \addr_calc/iir_write_addr[11] ,
         \addr_calc/iir_write_addr[10] , \addr_calc/iir_write_addr[9] ,
         \addr_calc/iir_write_addr[8] , \addr_calc/iir_write_addr[7] ,
         \addr_calc/iir_write_addr[6] , \addr_calc/iir_write_addr[5] ,
         \addr_calc/iir_write_addr[4] , \addr_calc/iir_write_addr[3] ,
         \addr_calc/iir_write_addr[2] , \addr_calc/iir_write_addr[1] ,
         \addr_calc/iir_write_addr[0] , \addr_calc/iir_read_addr[31] ,
         \addr_calc/iir_read_addr[30] , \addr_calc/iir_read_addr[29] ,
         \addr_calc/iir_read_addr[28] , \addr_calc/iir_read_addr[27] ,
         \addr_calc/iir_read_addr[26] , \addr_calc/iir_read_addr[25] ,
         \addr_calc/iir_read_addr[24] , \addr_calc/iir_read_addr[23] ,
         \addr_calc/iir_read_addr[22] , \addr_calc/iir_read_addr[21] ,
         \addr_calc/iir_read_addr[20] , \addr_calc/iir_read_addr[19] ,
         \addr_calc/iir_read_addr[18] , \addr_calc/iir_read_addr[17] ,
         \addr_calc/iir_read_addr[16] , \addr_calc/iir_read_addr[15] ,
         \addr_calc/iir_read_addr[14] , \addr_calc/iir_read_addr[13] ,
         \addr_calc/iir_read_addr[12] , \addr_calc/iir_read_addr[11] ,
         \addr_calc/iir_read_addr[10] , \addr_calc/iir_read_addr[9] ,
         \addr_calc/iir_read_addr[8] , \addr_calc/iir_read_addr[7] ,
         \addr_calc/iir_read_addr[6] , \addr_calc/iir_read_addr[5] ,
         \addr_calc/iir_read_addr[4] , \addr_calc/iir_read_addr[3] ,
         \addr_calc/iir_read_addr[2] , \addr_calc/iir_read_addr[1] ,
         \addr_calc/iir_read_addr[0] , \addr_calc/fir_write_addr[31] ,
         \addr_calc/fir_write_addr[30] , \addr_calc/fir_write_addr[29] ,
         \addr_calc/fir_write_addr[28] , \addr_calc/fir_write_addr[27] ,
         \addr_calc/fir_write_addr[26] , \addr_calc/fir_write_addr[25] ,
         \addr_calc/fir_write_addr[24] , \addr_calc/fir_write_addr[23] ,
         \addr_calc/fir_write_addr[22] , \addr_calc/fir_write_addr[21] ,
         \addr_calc/fir_write_addr[20] , \addr_calc/fir_write_addr[19] ,
         \addr_calc/fir_write_addr[18] , \addr_calc/fir_write_addr[17] ,
         \addr_calc/fir_write_addr[16] , \addr_calc/fir_write_addr[15] ,
         \addr_calc/fir_write_addr[14] , \addr_calc/fir_write_addr[13] ,
         \addr_calc/fir_write_addr[12] , \addr_calc/fir_write_addr[11] ,
         \addr_calc/fir_write_addr[10] , \addr_calc/fir_write_addr[9] ,
         \addr_calc/fir_write_addr[8] , \addr_calc/fir_write_addr[7] ,
         \addr_calc/fir_write_addr[6] , \addr_calc/fir_write_addr[5] ,
         \addr_calc/fir_write_addr[4] , \addr_calc/fir_write_addr[3] ,
         \addr_calc/fir_write_addr[2] , \addr_calc/fir_write_addr[1] ,
         \addr_calc/fir_write_addr[0] , \addr_calc/fir_read_addr[31] ,
         \addr_calc/fir_read_addr[30] , \addr_calc/fir_read_addr[29] ,
         \addr_calc/fir_read_addr[28] , \addr_calc/fir_read_addr[27] ,
         \addr_calc/fir_read_addr[26] , \addr_calc/fir_read_addr[25] ,
         \addr_calc/fir_read_addr[24] , \addr_calc/fir_read_addr[23] ,
         \addr_calc/fir_read_addr[22] , \addr_calc/fir_read_addr[21] ,
         \addr_calc/fir_read_addr[20] , \addr_calc/fir_read_addr[19] ,
         \addr_calc/fir_read_addr[18] , \addr_calc/fir_read_addr[17] ,
         \addr_calc/fir_read_addr[16] , \addr_calc/fir_read_addr[15] ,
         \addr_calc/fir_read_addr[14] , \addr_calc/fir_read_addr[13] ,
         \addr_calc/fir_read_addr[12] , \addr_calc/fir_read_addr[11] ,
         \addr_calc/fir_read_addr[10] , \addr_calc/fir_read_addr[9] ,
         \addr_calc/fir_read_addr[8] , \addr_calc/fir_read_addr[7] ,
         \addr_calc/fir_read_addr[6] , \addr_calc/fir_read_addr[5] ,
         \addr_calc/fir_read_addr[4] , \addr_calc/fir_read_addr[3] ,
         \addr_calc/fir_read_addr[2] , \addr_calc/fir_read_addr[1] ,
         \addr_calc/fir_read_addr[0] , \addr_calc/fft_write_addr[31] ,
         \addr_calc/fft_write_addr[30] , \addr_calc/fft_write_addr[29] ,
         \addr_calc/fft_write_addr[28] , \addr_calc/fft_write_addr[27] ,
         \addr_calc/fft_write_addr[26] , \addr_calc/fft_write_addr[25] ,
         \addr_calc/fft_write_addr[24] , \addr_calc/fft_write_addr[23] ,
         \addr_calc/fft_write_addr[22] , \addr_calc/fft_write_addr[21] ,
         \addr_calc/fft_write_addr[20] , \addr_calc/fft_write_addr[19] ,
         \addr_calc/fft_write_addr[18] , \addr_calc/fft_write_addr[17] ,
         \addr_calc/fft_write_addr[16] , \addr_calc/fft_write_addr[15] ,
         \addr_calc/fft_write_addr[14] , \addr_calc/fft_write_addr[13] ,
         \addr_calc/fft_write_addr[12] , \addr_calc/fft_write_addr[11] ,
         \addr_calc/fft_write_addr[10] , \addr_calc/fft_write_addr[9] ,
         \addr_calc/fft_write_addr[8] , \addr_calc/fft_write_addr[7] ,
         \addr_calc/fft_write_addr[6] , \addr_calc/fft_write_addr[5] ,
         \addr_calc/fft_write_addr[4] , \addr_calc/fft_write_addr[3] ,
         \addr_calc/fft_write_addr[2] , \addr_calc/fft_write_addr[1] ,
         \addr_calc/fft_write_addr[0] , \addr_calc/fft_read_addr[31] ,
         \addr_calc/fft_read_addr[30] , \addr_calc/fft_read_addr[29] ,
         \addr_calc/fft_read_addr[28] , \addr_calc/fft_read_addr[27] ,
         \addr_calc/fft_read_addr[26] , \addr_calc/fft_read_addr[25] ,
         \addr_calc/fft_read_addr[24] , \addr_calc/fft_read_addr[23] ,
         \addr_calc/fft_read_addr[22] , \addr_calc/fft_read_addr[21] ,
         \addr_calc/fft_read_addr[20] , \addr_calc/fft_read_addr[19] ,
         \addr_calc/fft_read_addr[18] , \addr_calc/fft_read_addr[17] ,
         \addr_calc/fft_read_addr[16] , \addr_calc/fft_read_addr[15] ,
         \addr_calc/fft_read_addr[14] , \addr_calc/fft_read_addr[13] ,
         \addr_calc/fft_read_addr[12] , \addr_calc/fft_read_addr[11] ,
         \addr_calc/fft_read_addr[10] , \addr_calc/fft_read_addr[9] ,
         \addr_calc/fft_read_addr[8] , \addr_calc/fft_read_addr[7] ,
         \addr_calc/fft_read_addr[6] , \addr_calc/fft_read_addr[5] ,
         \addr_calc/fft_read_addr[4] , \addr_calc/fft_read_addr[3] ,
         \addr_calc/fft_read_addr[2] , \addr_calc/fft_read_addr[1] ,
         \addr_calc/fft_read_addr[0] , \addr_calc/N191 , \addr_calc/N159 ,
         \addr_calc/N99 , \addr_calc/N95 , \addr_calc/N63 , \addr_calc/N9 ,
         \data_cntl/N267 , \data_cntl/N266 , \data_cntl/N265 ,
         \data_cntl/N264 , \data_cntl/N263 , \data_cntl/N262 ,
         \data_cntl/N261 , \data_cntl/N260 , \data_cntl/N259 ,
         \data_cntl/N258 , \data_cntl/N257 , \data_cntl/N256 ,
         \data_cntl/N255 , \data_cntl/N254 , \data_cntl/N253 ,
         \data_cntl/N252 , \data_cntl/N251 , \data_cntl/N250 ,
         \data_cntl/N191 , \data_cntl/N159 , \data_cntl/N99 , \data_cntl/N95 ,
         \data_cntl/N63 , \data_cntl/N9 , \addr_calc/fft_read_calc/count[31] ,
         \addr_calc/fft_read_calc/count[30] ,
         \addr_calc/fft_read_calc/count[29] ,
         \addr_calc/fft_read_calc/count[28] ,
         \addr_calc/fft_read_calc/count[27] ,
         \addr_calc/fft_read_calc/count[26] ,
         \addr_calc/fft_read_calc/count[25] ,
         \addr_calc/fft_read_calc/count[24] ,
         \addr_calc/fft_read_calc/count[23] ,
         \addr_calc/fft_read_calc/count[22] ,
         \addr_calc/fft_read_calc/count[21] ,
         \addr_calc/fft_read_calc/count[20] ,
         \addr_calc/fft_read_calc/count[19] ,
         \addr_calc/fft_read_calc/count[18] ,
         \addr_calc/fft_read_calc/count[17] ,
         \addr_calc/fft_read_calc/count[16] ,
         \addr_calc/fft_read_calc/count[15] ,
         \addr_calc/fft_read_calc/count[14] ,
         \addr_calc/fft_read_calc/count[13] ,
         \addr_calc/fft_read_calc/count[12] ,
         \addr_calc/fft_read_calc/count[11] ,
         \addr_calc/fft_read_calc/count[10] ,
         \addr_calc/fft_read_calc/count[9] ,
         \addr_calc/fft_read_calc/count[8] ,
         \addr_calc/fft_read_calc/count[7] ,
         \addr_calc/fft_read_calc/count[6] ,
         \addr_calc/fft_read_calc/count[5] ,
         \addr_calc/fft_read_calc/count[4] ,
         \addr_calc/fft_read_calc/count[3] ,
         \addr_calc/fft_read_calc/count[2] ,
         \addr_calc/fft_read_calc/count[1] ,
         \addr_calc/fft_read_calc/count[0] ,
         \addr_calc/fft_write_calc/count[31] ,
         \addr_calc/fft_write_calc/count[30] ,
         \addr_calc/fft_write_calc/count[29] ,
         \addr_calc/fft_write_calc/count[28] ,
         \addr_calc/fft_write_calc/count[27] ,
         \addr_calc/fft_write_calc/count[26] ,
         \addr_calc/fft_write_calc/count[25] ,
         \addr_calc/fft_write_calc/count[24] ,
         \addr_calc/fft_write_calc/count[23] ,
         \addr_calc/fft_write_calc/count[22] ,
         \addr_calc/fft_write_calc/count[21] ,
         \addr_calc/fft_write_calc/count[20] ,
         \addr_calc/fft_write_calc/count[19] ,
         \addr_calc/fft_write_calc/count[18] ,
         \addr_calc/fft_write_calc/count[17] ,
         \addr_calc/fft_write_calc/count[16] ,
         \addr_calc/fft_write_calc/count[15] ,
         \addr_calc/fft_write_calc/count[14] ,
         \addr_calc/fft_write_calc/count[13] ,
         \addr_calc/fft_write_calc/count[12] ,
         \addr_calc/fft_write_calc/count[11] ,
         \addr_calc/fft_write_calc/count[10] ,
         \addr_calc/fft_write_calc/count[9] ,
         \addr_calc/fft_write_calc/count[8] ,
         \addr_calc/fft_write_calc/count[7] ,
         \addr_calc/fft_write_calc/count[6] ,
         \addr_calc/fft_write_calc/count[5] ,
         \addr_calc/fft_write_calc/count[4] ,
         \addr_calc/fft_write_calc/count[3] ,
         \addr_calc/fft_write_calc/count[2] ,
         \addr_calc/fft_write_calc/count[1] ,
         \addr_calc/fft_write_calc/count[0] ,
         \addr_calc/fir_read_calc/count[31] ,
         \addr_calc/fir_read_calc/count[30] ,
         \addr_calc/fir_read_calc/count[29] ,
         \addr_calc/fir_read_calc/count[28] ,
         \addr_calc/fir_read_calc/count[27] ,
         \addr_calc/fir_read_calc/count[26] ,
         \addr_calc/fir_read_calc/count[25] ,
         \addr_calc/fir_read_calc/count[24] ,
         \addr_calc/fir_read_calc/count[23] ,
         \addr_calc/fir_read_calc/count[22] ,
         \addr_calc/fir_read_calc/count[21] ,
         \addr_calc/fir_read_calc/count[20] ,
         \addr_calc/fir_read_calc/count[19] ,
         \addr_calc/fir_read_calc/count[18] ,
         \addr_calc/fir_read_calc/count[17] ,
         \addr_calc/fir_read_calc/count[16] ,
         \addr_calc/fir_read_calc/count[15] ,
         \addr_calc/fir_read_calc/count[14] ,
         \addr_calc/fir_read_calc/count[13] ,
         \addr_calc/fir_read_calc/count[12] ,
         \addr_calc/fir_read_calc/count[11] ,
         \addr_calc/fir_read_calc/count[10] ,
         \addr_calc/fir_read_calc/count[9] ,
         \addr_calc/fir_read_calc/count[8] ,
         \addr_calc/fir_read_calc/count[7] ,
         \addr_calc/fir_read_calc/count[6] ,
         \addr_calc/fir_read_calc/count[5] ,
         \addr_calc/fir_read_calc/count[4] ,
         \addr_calc/fir_read_calc/count[3] ,
         \addr_calc/fir_read_calc/count[2] ,
         \addr_calc/fir_read_calc/count[1] ,
         \addr_calc/fir_read_calc/count[0] ,
         \addr_calc/fir_write_calc/count[31] ,
         \addr_calc/fir_write_calc/count[30] ,
         \addr_calc/fir_write_calc/count[29] ,
         \addr_calc/fir_write_calc/count[28] ,
         \addr_calc/fir_write_calc/count[27] ,
         \addr_calc/fir_write_calc/count[26] ,
         \addr_calc/fir_write_calc/count[25] ,
         \addr_calc/fir_write_calc/count[24] ,
         \addr_calc/fir_write_calc/count[23] ,
         \addr_calc/fir_write_calc/count[22] ,
         \addr_calc/fir_write_calc/count[21] ,
         \addr_calc/fir_write_calc/count[20] ,
         \addr_calc/fir_write_calc/count[19] ,
         \addr_calc/fir_write_calc/count[18] ,
         \addr_calc/fir_write_calc/count[17] ,
         \addr_calc/fir_write_calc/count[16] ,
         \addr_calc/fir_write_calc/count[15] ,
         \addr_calc/fir_write_calc/count[14] ,
         \addr_calc/fir_write_calc/count[13] ,
         \addr_calc/fir_write_calc/count[12] ,
         \addr_calc/fir_write_calc/count[11] ,
         \addr_calc/fir_write_calc/count[10] ,
         \addr_calc/fir_write_calc/count[9] ,
         \addr_calc/fir_write_calc/count[8] ,
         \addr_calc/fir_write_calc/count[7] ,
         \addr_calc/fir_write_calc/count[6] ,
         \addr_calc/fir_write_calc/count[5] ,
         \addr_calc/fir_write_calc/count[4] ,
         \addr_calc/fir_write_calc/count[3] ,
         \addr_calc/fir_write_calc/count[2] ,
         \addr_calc/fir_write_calc/count[1] ,
         \addr_calc/fir_write_calc/count[0] ,
         \addr_calc/iir_read_calc/count[31] ,
         \addr_calc/iir_read_calc/count[30] ,
         \addr_calc/iir_read_calc/count[29] ,
         \addr_calc/iir_read_calc/count[28] ,
         \addr_calc/iir_read_calc/count[27] ,
         \addr_calc/iir_read_calc/count[26] ,
         \addr_calc/iir_read_calc/count[25] ,
         \addr_calc/iir_read_calc/count[24] ,
         \addr_calc/iir_read_calc/count[23] ,
         \addr_calc/iir_read_calc/count[22] ,
         \addr_calc/iir_read_calc/count[21] ,
         \addr_calc/iir_read_calc/count[20] ,
         \addr_calc/iir_read_calc/count[19] ,
         \addr_calc/iir_read_calc/count[18] ,
         \addr_calc/iir_read_calc/count[17] ,
         \addr_calc/iir_read_calc/count[16] ,
         \addr_calc/iir_read_calc/count[15] ,
         \addr_calc/iir_read_calc/count[14] ,
         \addr_calc/iir_read_calc/count[13] ,
         \addr_calc/iir_read_calc/count[12] ,
         \addr_calc/iir_read_calc/count[11] ,
         \addr_calc/iir_read_calc/count[10] ,
         \addr_calc/iir_read_calc/count[9] ,
         \addr_calc/iir_read_calc/count[8] ,
         \addr_calc/iir_read_calc/count[7] ,
         \addr_calc/iir_read_calc/count[6] ,
         \addr_calc/iir_read_calc/count[5] ,
         \addr_calc/iir_read_calc/count[4] ,
         \addr_calc/iir_read_calc/count[3] ,
         \addr_calc/iir_read_calc/count[2] ,
         \addr_calc/iir_read_calc/count[1] ,
         \addr_calc/iir_read_calc/count[0] ,
         \addr_calc/iir_write_calc/count[31] ,
         \addr_calc/iir_write_calc/count[30] ,
         \addr_calc/iir_write_calc/count[29] ,
         \addr_calc/iir_write_calc/count[28] ,
         \addr_calc/iir_write_calc/count[27] ,
         \addr_calc/iir_write_calc/count[26] ,
         \addr_calc/iir_write_calc/count[25] ,
         \addr_calc/iir_write_calc/count[24] ,
         \addr_calc/iir_write_calc/count[23] ,
         \addr_calc/iir_write_calc/count[22] ,
         \addr_calc/iir_write_calc/count[21] ,
         \addr_calc/iir_write_calc/count[20] ,
         \addr_calc/iir_write_calc/count[19] ,
         \addr_calc/iir_write_calc/count[18] ,
         \addr_calc/iir_write_calc/count[17] ,
         \addr_calc/iir_write_calc/count[16] ,
         \addr_calc/iir_write_calc/count[15] ,
         \addr_calc/iir_write_calc/count[14] ,
         \addr_calc/iir_write_calc/count[13] ,
         \addr_calc/iir_write_calc/count[12] ,
         \addr_calc/iir_write_calc/count[11] ,
         \addr_calc/iir_write_calc/count[10] ,
         \addr_calc/iir_write_calc/count[9] ,
         \addr_calc/iir_write_calc/count[8] ,
         \addr_calc/iir_write_calc/count[7] ,
         \addr_calc/iir_write_calc/count[6] ,
         \addr_calc/iir_write_calc/count[5] ,
         \addr_calc/iir_write_calc/count[4] ,
         \addr_calc/iir_write_calc/count[3] ,
         \addr_calc/iir_write_calc/count[2] ,
         \addr_calc/iir_write_calc/count[1] ,
         \addr_calc/iir_write_calc/count[0] ,
         \addr_calc/fft_read_calc/counter/N73 ,
         \addr_calc/fft_read_calc/counter/N72 ,
         \addr_calc/fft_read_calc/counter/N71 ,
         \addr_calc/fft_read_calc/counter/N70 ,
         \addr_calc/fft_read_calc/counter/N68 ,
         \addr_calc/fft_read_calc/counter/N67 ,
         \addr_calc/fft_read_calc/counter/N66 ,
         \addr_calc/fft_read_calc/counter/N65 ,
         \addr_calc/fft_read_calc/counter/N63 ,
         \addr_calc/fft_read_calc/counter/N62 ,
         \addr_calc/fft_read_calc/counter/N58 ,
         \addr_calc/fft_read_calc/counter/N57 ,
         \addr_calc/fft_read_calc/counter/N56 ,
         \addr_calc/fft_read_calc/counter/N55 ,
         \addr_calc/fft_read_calc/counter/N53 ,
         \addr_calc/fft_read_calc/counter/N52 ,
         \addr_calc/fft_read_calc/counter/N51 ,
         \addr_calc/fft_read_calc/counter/N50 ,
         \addr_calc/fft_read_calc/counter/N48 ,
         \addr_calc/fft_read_calc/counter/N46 ,
         \addr_calc/fft_read_calc/counter/N45 ,
         \addr_calc/fft_read_calc/counter/N44 ,
         \addr_calc/fft_read_calc/counter/N38 ,
         \addr_calc/fft_write_calc/counter/N74 ,
         \addr_calc/fft_write_calc/counter/N73 ,
         \addr_calc/fft_write_calc/counter/N72 ,
         \addr_calc/fft_write_calc/counter/N71 ,
         \addr_calc/fft_write_calc/counter/N68 ,
         \addr_calc/fft_write_calc/counter/N66 ,
         \addr_calc/fft_write_calc/counter/N64 ,
         \addr_calc/fft_write_calc/counter/N62 ,
         \addr_calc/fft_write_calc/counter/N60 ,
         \addr_calc/fft_write_calc/counter/N59 ,
         \addr_calc/fft_write_calc/counter/N58 ,
         \addr_calc/fft_write_calc/counter/N57 ,
         \addr_calc/fft_write_calc/counter/N56 ,
         \addr_calc/fft_write_calc/counter/N55 ,
         \addr_calc/fft_write_calc/counter/N53 ,
         \addr_calc/fft_write_calc/counter/N52 ,
         \addr_calc/fft_write_calc/counter/N51 ,
         \addr_calc/fft_write_calc/counter/N50 ,
         \addr_calc/fft_write_calc/counter/N47 ,
         \addr_calc/fft_write_calc/counter/N46 ,
         \addr_calc/fft_write_calc/counter/N43 ,
         \addr_calc/fft_write_calc/counter/N38 ,
         \addr_calc/fir_read_calc/counter/N73 ,
         \addr_calc/fir_read_calc/counter/N72 ,
         \addr_calc/fir_read_calc/counter/N71 ,
         \addr_calc/fir_read_calc/counter/N67 ,
         \addr_calc/fir_read_calc/counter/N66 ,
         \addr_calc/fir_read_calc/counter/N65 ,
         \addr_calc/fir_read_calc/counter/N64 ,
         \addr_calc/fir_read_calc/counter/N63 ,
         \addr_calc/fir_read_calc/counter/N62 ,
         \addr_calc/fir_read_calc/counter/N61 ,
         \addr_calc/fir_read_calc/counter/N60 ,
         \addr_calc/fir_read_calc/counter/N59 ,
         \addr_calc/fir_read_calc/counter/N57 ,
         \addr_calc/fir_read_calc/counter/N56 ,
         \addr_calc/fir_read_calc/counter/N55 ,
         \addr_calc/fir_read_calc/counter/N54 ,
         \addr_calc/fir_read_calc/counter/N53 ,
         \addr_calc/fir_read_calc/counter/N52 ,
         \addr_calc/fir_read_calc/counter/N51 ,
         \addr_calc/fir_read_calc/counter/N50 ,
         \addr_calc/fir_read_calc/counter/N49 ,
         \addr_calc/fir_read_calc/counter/N48 ,
         \addr_calc/fir_read_calc/counter/N47 ,
         \addr_calc/fir_read_calc/counter/N45 ,
         \addr_calc/fir_read_calc/counter/N44 ,
         \addr_calc/fir_read_calc/counter/N38 ,
         \addr_calc/fir_write_calc/counter/N74 ,
         \addr_calc/fir_write_calc/counter/N73 ,
         \addr_calc/fir_write_calc/counter/N72 ,
         \addr_calc/fir_write_calc/counter/N71 ,
         \addr_calc/fir_write_calc/counter/N70 ,
         \addr_calc/fir_write_calc/counter/N68 ,
         \addr_calc/fir_write_calc/counter/N67 ,
         \addr_calc/fir_write_calc/counter/N66 ,
         \addr_calc/fir_write_calc/counter/N65 ,
         \addr_calc/fir_write_calc/counter/N62 ,
         \addr_calc/fir_write_calc/counter/N61 ,
         \addr_calc/fir_write_calc/counter/N60 ,
         \addr_calc/fir_write_calc/counter/N59 ,
         \addr_calc/fir_write_calc/counter/N57 ,
         \addr_calc/fir_write_calc/counter/N56 ,
         \addr_calc/fir_write_calc/counter/N54 ,
         \addr_calc/fir_write_calc/counter/N52 ,
         \addr_calc/fir_write_calc/counter/N51 ,
         \addr_calc/fir_write_calc/counter/N49 ,
         \addr_calc/fir_write_calc/counter/N48 ,
         \addr_calc/fir_write_calc/counter/N46 ,
         \addr_calc/fir_write_calc/counter/N45 ,
         \addr_calc/fir_write_calc/counter/N43 ,
         \addr_calc/fir_write_calc/counter/N38 ,
         \addr_calc/iir_read_calc/counter/N74 ,
         \addr_calc/iir_read_calc/counter/N73 ,
         \addr_calc/iir_read_calc/counter/N72 ,
         \addr_calc/iir_read_calc/counter/N71 ,
         \addr_calc/iir_read_calc/counter/N68 ,
         \addr_calc/iir_read_calc/counter/N67 ,
         \addr_calc/iir_read_calc/counter/N63 ,
         \addr_calc/iir_read_calc/counter/N62 ,
         \addr_calc/iir_read_calc/counter/N61 ,
         \addr_calc/iir_read_calc/counter/N60 ,
         \addr_calc/iir_read_calc/counter/N59 ,
         \addr_calc/iir_read_calc/counter/N58 ,
         \addr_calc/iir_read_calc/counter/N57 ,
         \addr_calc/iir_read_calc/counter/N55 ,
         \addr_calc/iir_read_calc/counter/N54 ,
         \addr_calc/iir_read_calc/counter/N53 ,
         \addr_calc/iir_read_calc/counter/N52 ,
         \addr_calc/iir_read_calc/counter/N51 ,
         \addr_calc/iir_read_calc/counter/N50 ,
         \addr_calc/iir_read_calc/counter/N48 ,
         \addr_calc/iir_read_calc/counter/N46 ,
         \addr_calc/iir_read_calc/counter/N45 ,
         \addr_calc/iir_read_calc/counter/N44 ,
         \addr_calc/iir_write_calc/counter/N74 ,
         \addr_calc/iir_write_calc/counter/N73 ,
         \addr_calc/iir_write_calc/counter/N72 ,
         \addr_calc/iir_write_calc/counter/N71 ,
         \addr_calc/iir_write_calc/counter/N70 ,
         \addr_calc/iir_write_calc/counter/N69 ,
         \addr_calc/iir_write_calc/counter/N68 ,
         \addr_calc/iir_write_calc/counter/N67 ,
         \addr_calc/iir_write_calc/counter/N66 ,
         \addr_calc/iir_write_calc/counter/N65 ,
         \addr_calc/iir_write_calc/counter/N62 ,
         \addr_calc/iir_write_calc/counter/N60 ,
         \addr_calc/iir_write_calc/counter/N57 ,
         \addr_calc/iir_write_calc/counter/N56 ,
         \addr_calc/iir_write_calc/counter/N55 ,
         \addr_calc/iir_write_calc/counter/N54 ,
         \addr_calc/iir_write_calc/counter/N53 ,
         \addr_calc/iir_write_calc/counter/N52 ,
         \addr_calc/iir_write_calc/counter/N51 ,
         \addr_calc/iir_write_calc/counter/N50 ,
         \addr_calc/iir_write_calc/counter/N49 ,
         \addr_calc/iir_write_calc/counter/N48 ,
         \addr_calc/iir_write_calc/counter/N47 ,
         \addr_calc/iir_write_calc/counter/N46 ,
         \addr_calc/iir_write_calc/counter/N45 ,
         \addr_calc/iir_write_calc/counter/N44 , n3, n67, n131, n195, n259,
         n323, n387, n451, n515, n579, n643, n707, n783, n785, n787, n790,
         n791, n792, n793, n795, n796, n797, n798, n801, n802, n810, n811,
         n812, n813, n814, n815, n816, n817, n828, n829, n830, n831, n832,
         n833, n842, n843, n844, n845, n846, n847, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, \add_x_19_4/n222 , \add_x_19_4/n221 , \add_x_19_4/n219 ,
         \add_x_19_4/n217 , \add_x_19_4/n213 , \add_x_19_4/n212 ,
         \add_x_19_4/n207 , \add_x_19_4/n206 , \add_x_19_4/n204 ,
         \add_x_19_4/n202 , \add_x_19_4/n199 , \add_x_19_4/n196 ,
         \add_x_19_4/n191 , \add_x_19_4/n189 , \add_x_19_4/n188 ,
         \add_x_19_4/n187 , \add_x_19_4/n186 , \add_x_19_4/n185 ,
         \add_x_19_4/n184 , \add_x_19_4/n182 , \add_x_19_4/n181 ,
         \add_x_19_4/n178 , \add_x_19_4/n177 , \add_x_19_4/n176 ,
         \add_x_19_4/n175 , \add_x_19_4/n171 , \add_x_19_4/n170 ,
         \add_x_19_4/n169 , \add_x_19_4/n168 , \add_x_19_4/n167 ,
         \add_x_19_4/n166 , \add_x_19_4/n165 , \add_x_19_4/n163 ,
         \add_x_19_4/n162 , \add_x_19_4/n160 , \add_x_19_4/n157 ,
         \add_x_19_4/n156 , \add_x_19_4/n155 , \add_x_19_4/n154 ,
         \add_x_19_4/n152 , \add_x_19_4/n151 , \add_x_19_4/n150 ,
         \add_x_19_4/n149 , \add_x_19_4/n148 , \add_x_19_4/n147 ,
         \add_x_19_4/n146 , \add_x_19_4/n145 , \add_x_19_4/n144 ,
         \add_x_19_4/n143 , \add_x_19_4/n141 , \add_x_19_4/n140 ,
         \add_x_19_4/n139 , \add_x_19_4/n138 , \add_x_19_4/n137 ,
         \add_x_19_4/n136 , \add_x_19_4/n135 , \add_x_19_4/n134 ,
         \add_x_19_4/n133 , \add_x_19_4/n132 , \add_x_19_4/n131 ,
         \add_x_19_4/n130 , \add_x_19_4/n129 , \add_x_19_4/n128 ,
         \add_x_19_4/n127 , \add_x_19_4/n126 , \add_x_19_4/n125 ,
         \add_x_19_4/n124 , \add_x_19_4/n123 , \add_x_19_4/n121 ,
         \add_x_19_4/n120 , \add_x_19_4/n112 , \add_x_19_4/n111 ,
         \add_x_19_4/n110 , \add_x_19_4/n109 , \add_x_19_4/n107 ,
         \add_x_19_4/n106 , \add_x_19_4/n105 , \add_x_19_4/n104 ,
         \add_x_19_4/n103 , \add_x_19_4/n102 , \add_x_19_4/n101 ,
         \add_x_19_4/n100 , \add_x_19_4/n99 , \add_x_19_4/n98 ,
         \add_x_19_4/n97 , \add_x_19_4/n96 , \add_x_19_4/n95 ,
         \add_x_19_4/n94 , \add_x_19_4/n93 , \add_x_19_4/n91 ,
         \add_x_19_4/n90 , \add_x_19_4/n89 , \add_x_19_4/n88 ,
         \add_x_19_4/n87 , \add_x_19_4/n86 , \add_x_19_4/n85 ,
         \add_x_19_4/n84 , \add_x_19_4/n82 , \add_x_19_4/n81 ,
         \add_x_19_4/n79 , \add_x_19_4/n78 , \add_x_19_4/n77 ,
         \add_x_19_4/n76 , \add_x_19_4/n75 , \add_x_19_4/n74 ,
         \add_x_19_4/n73 , \add_x_19_4/n72 , \add_x_19_4/n69 ,
         \add_x_19_4/n67 , \add_x_19_4/n66 , \add_x_19_4/n64 ,
         \add_x_19_4/n63 , \add_x_19_4/n62 , \add_x_19_4/n61 ,
         \add_x_19_4/n60 , \add_x_19_4/n59 , \add_x_19_4/n58 ,
         \add_x_19_4/n57 , \add_x_19_4/n56 , \add_x_19_4/n55 ,
         \add_x_19_4/n54 , \add_x_19_4/n53 , \add_x_19_4/n52 ,
         \add_x_19_4/n51 , \add_x_19_4/n49 , \add_x_19_4/n48 ,
         \add_x_19_4/n46 , \add_x_19_4/n43 , \add_x_19_4/n42 ,
         \add_x_19_4/n37 , \add_x_19_4/n36 , \add_x_19_4/n31 ,
         \add_x_19_4/n30 , \add_x_19_4/n28 , \add_x_19_4/n26 ,
         \add_x_19_4/n22 , \add_x_19_4/n21 , \add_x_19_4/n19 ,
         \add_x_19_4/n15 , \add_x_19_4/n13 , \add_x_19_4/n11 , \add_x_19_4/n5 ,
         \add_x_19_4/n3 , \add_x_19_2/n219 , \add_x_19_2/n216 ,
         \add_x_19_2/n215 , \add_x_19_2/n213 , \add_x_19_2/n212 ,
         \add_x_19_2/n210 , \add_x_19_2/n208 , \add_x_19_2/n207 ,
         \add_x_19_2/n206 , \add_x_19_2/n204 , \add_x_19_2/n191 ,
         \add_x_19_2/n189 , \add_x_19_2/n188 , \add_x_19_2/n187 ,
         \add_x_19_2/n186 , \add_x_19_2/n185 , \add_x_19_2/n184 ,
         \add_x_19_2/n182 , \add_x_19_2/n181 , \add_x_19_2/n178 ,
         \add_x_19_2/n177 , \add_x_19_2/n176 , \add_x_19_2/n175 ,
         \add_x_19_2/n171 , \add_x_19_2/n170 , \add_x_19_2/n169 ,
         \add_x_19_2/n168 , \add_x_19_2/n167 , \add_x_19_2/n166 ,
         \add_x_19_2/n165 , \add_x_19_2/n164 , \add_x_19_2/n163 ,
         \add_x_19_2/n156 , \add_x_19_2/n155 , \add_x_19_2/n154 ,
         \add_x_19_2/n152 , \add_x_19_2/n151 , \add_x_19_2/n150 ,
         \add_x_19_2/n149 , \add_x_19_2/n148 , \add_x_19_2/n147 ,
         \add_x_19_2/n146 , \add_x_19_2/n144 , \add_x_19_2/n143 ,
         \add_x_19_2/n140 , \add_x_19_2/n139 , \add_x_19_2/n137 ,
         \add_x_19_2/n135 , \add_x_19_2/n134 , \add_x_19_2/n133 ,
         \add_x_19_2/n132 , \add_x_19_2/n131 , \add_x_19_2/n130 ,
         \add_x_19_2/n129 , \add_x_19_2/n128 , \add_x_19_2/n127 ,
         \add_x_19_2/n126 , \add_x_19_2/n125 , \add_x_19_2/n124 ,
         \add_x_19_2/n123 , \add_x_19_2/n122 , \add_x_19_2/n121 ,
         \add_x_19_2/n120 , \add_x_19_2/n118 , \add_x_19_2/n116 ,
         \add_x_19_2/n112 , \add_x_19_2/n111 , \add_x_19_2/n110 ,
         \add_x_19_2/n109 , \add_x_19_2/n107 , \add_x_19_2/n106 ,
         \add_x_19_2/n105 , \add_x_19_2/n104 , \add_x_19_2/n103 ,
         \add_x_19_2/n102 , \add_x_19_2/n101 , \add_x_19_2/n100 ,
         \add_x_19_2/n99 , \add_x_19_2/n98 , \add_x_19_2/n97 ,
         \add_x_19_2/n96 , \add_x_19_2/n95 , \add_x_19_2/n94 ,
         \add_x_19_2/n93 , \add_x_19_2/n92 , \add_x_19_2/n91 ,
         \add_x_19_2/n90 , \add_x_19_2/n89 , \add_x_19_2/n87 ,
         \add_x_19_2/n86 , \add_x_19_2/n85 , \add_x_19_2/n84 ,
         \add_x_19_2/n83 , \add_x_19_2/n82 , \add_x_19_2/n81 ,
         \add_x_19_2/n79 , \add_x_19_2/n78 , \add_x_19_2/n76 ,
         \add_x_19_2/n74 , \add_x_19_2/n73 , \add_x_19_2/n72 ,
         \add_x_19_2/n69 , \add_x_19_2/n68 , \add_x_19_2/n67 ,
         \add_x_19_2/n66 , \add_x_19_2/n64 , \add_x_19_2/n63 ,
         \add_x_19_2/n62 , \add_x_19_2/n61 , \add_x_19_2/n60 ,
         \add_x_19_2/n59 , \add_x_19_2/n58 , \add_x_19_2/n56 ,
         \add_x_19_2/n55 , \add_x_19_2/n54 , \add_x_19_2/n53 ,
         \add_x_19_2/n52 , \add_x_19_2/n51 , \add_x_19_2/n49 ,
         \add_x_19_2/n48 , \add_x_19_2/n46 , \add_x_19_2/n42 ,
         \add_x_19_2/n37 , \add_x_19_2/n36 , \add_x_19_2/n28 ,
         \add_x_19_2/n25 , \add_x_19_2/n24 , \add_x_19_2/n19 ,
         \add_x_19_2/n17 , \add_x_19_2/n15 , \add_x_19_1/n219 ,
         \add_x_19_1/n218 , \add_x_19_1/n213 , \add_x_19_1/n212 ,
         \add_x_19_1/n210 , \add_x_19_1/n208 , \add_x_19_1/n207 ,
         \add_x_19_1/n202 , \add_x_19_1/n198 , \add_x_19_1/n195 ,
         \add_x_19_1/n191 , \add_x_19_1/n189 , \add_x_19_1/n188 ,
         \add_x_19_1/n187 , \add_x_19_1/n186 , \add_x_19_1/n185 ,
         \add_x_19_1/n184 , \add_x_19_1/n182 , \add_x_19_1/n181 ,
         \add_x_19_1/n178 , \add_x_19_1/n177 , \add_x_19_1/n176 ,
         \add_x_19_1/n175 , \add_x_19_1/n174 , \add_x_19_1/n172 ,
         \add_x_19_1/n168 , \add_x_19_1/n167 , \add_x_19_1/n166 ,
         \add_x_19_1/n165 , \add_x_19_1/n163 , \add_x_19_1/n162 ,
         \add_x_19_1/n160 , \add_x_19_1/n156 , \add_x_19_1/n155 ,
         \add_x_19_1/n154 , \add_x_19_1/n152 , \add_x_19_1/n151 ,
         \add_x_19_1/n150 , \add_x_19_1/n149 , \add_x_19_1/n148 ,
         \add_x_19_1/n147 , \add_x_19_1/n146 , \add_x_19_1/n145 ,
         \add_x_19_1/n144 , \add_x_19_1/n143 , \add_x_19_1/n141 ,
         \add_x_19_1/n140 , \add_x_19_1/n139 , \add_x_19_1/n137 ,
         \add_x_19_1/n136 , \add_x_19_1/n135 , \add_x_19_1/n134 ,
         \add_x_19_1/n133 , \add_x_19_1/n132 , \add_x_19_1/n131 ,
         \add_x_19_1/n130 , \add_x_19_1/n129 , \add_x_19_1/n128 ,
         \add_x_19_1/n127 , \add_x_19_1/n126 , \add_x_19_1/n125 ,
         \add_x_19_1/n124 , \add_x_19_1/n123 , \add_x_19_1/n122 ,
         \add_x_19_1/n121 , \add_x_19_1/n120 , \add_x_19_1/n118 ,
         \add_x_19_1/n116 , \add_x_19_1/n112 , \add_x_19_1/n111 ,
         \add_x_19_1/n110 , \add_x_19_1/n109 , \add_x_19_1/n106 ,
         \add_x_19_1/n105 , \add_x_19_1/n104 , \add_x_19_1/n103 ,
         \add_x_19_1/n102 , \add_x_19_1/n101 , \add_x_19_1/n100 ,
         \add_x_19_1/n98 , \add_x_19_1/n97 , \add_x_19_1/n96 ,
         \add_x_19_1/n95 , \add_x_19_1/n94 , \add_x_19_1/n93 ,
         \add_x_19_1/n91 , \add_x_19_1/n90 , \add_x_19_1/n89 ,
         \add_x_19_1/n88 , \add_x_19_1/n87 , \add_x_19_1/n86 ,
         \add_x_19_1/n85 , \add_x_19_1/n84 , \add_x_19_1/n82 ,
         \add_x_19_1/n81 , \add_x_19_1/n79 , \add_x_19_1/n78 ,
         \add_x_19_1/n77 , \add_x_19_1/n76 , \add_x_19_1/n75 ,
         \add_x_19_1/n74 , \add_x_19_1/n73 , \add_x_19_1/n72 ,
         \add_x_19_1/n69 , \add_x_19_1/n68 , \add_x_19_1/n67 ,
         \add_x_19_1/n66 , \add_x_19_1/n65 , \add_x_19_1/n64 ,
         \add_x_19_1/n63 , \add_x_19_1/n62 , \add_x_19_1/n61 ,
         \add_x_19_1/n60 , \add_x_19_1/n59 , \add_x_19_1/n58 ,
         \add_x_19_1/n56 , \add_x_19_1/n55 , \add_x_19_1/n54 ,
         \add_x_19_1/n53 , \add_x_19_1/n52 , \add_x_19_1/n51 ,
         \add_x_19_1/n50 , \add_x_19_1/n49 , \add_x_19_1/n48 ,
         \add_x_19_1/n47 , \add_x_19_1/n46 , \add_x_19_1/n45 ,
         \add_x_19_1/n44 , \add_x_19_1/n43 , \add_x_19_1/n42 ,
         \add_x_19_1/n38 , \add_x_19_1/n37 , \add_x_19_1/n36 ,
         \add_x_19_1/n28 , \add_x_19_1/n27 , \add_x_19_1/n21 ,
         \add_x_19_1/n19 , \add_x_19_1/n17 , \add_x_19_1/n11 , \add_x_19_1/n7 ,
         \add_x_19_1/n4 , \add_x_19_1/n3 , \add_x_19_3/n221 ,
         \add_x_19_3/n219 , \add_x_19_3/n218 , \add_x_19_3/n217 ,
         \add_x_19_3/n215 , \add_x_19_3/n213 , \add_x_19_3/n208 ,
         \add_x_19_3/n207 , \add_x_19_3/n204 , \add_x_19_3/n202 ,
         \add_x_19_3/n198 , \add_x_19_3/n195 , \add_x_19_3/n191 ,
         \add_x_19_3/n189 , \add_x_19_3/n188 , \add_x_19_3/n187 ,
         \add_x_19_3/n186 , \add_x_19_3/n185 , \add_x_19_3/n184 ,
         \add_x_19_3/n182 , \add_x_19_3/n181 , \add_x_19_3/n178 ,
         \add_x_19_3/n177 , \add_x_19_3/n176 , \add_x_19_3/n175 ,
         \add_x_19_3/n174 , \add_x_19_3/n172 , \add_x_19_3/n171 ,
         \add_x_19_3/n170 , \add_x_19_3/n169 , \add_x_19_3/n168 ,
         \add_x_19_3/n167 , \add_x_19_3/n166 , \add_x_19_3/n165 ,
         \add_x_19_3/n163 , \add_x_19_3/n162 , \add_x_19_3/n160 ,
         \add_x_19_3/n157 , \add_x_19_3/n156 , \add_x_19_3/n155 ,
         \add_x_19_3/n154 , \add_x_19_3/n152 , \add_x_19_3/n151 ,
         \add_x_19_3/n150 , \add_x_19_3/n149 , \add_x_19_3/n148 ,
         \add_x_19_3/n147 , \add_x_19_3/n146 , \add_x_19_3/n145 ,
         \add_x_19_3/n144 , \add_x_19_3/n140 , \add_x_19_3/n139 ,
         \add_x_19_3/n137 , \add_x_19_3/n136 , \add_x_19_3/n135 ,
         \add_x_19_3/n134 , \add_x_19_3/n133 , \add_x_19_3/n132 ,
         \add_x_19_3/n131 , \add_x_19_3/n129 , \add_x_19_3/n128 ,
         \add_x_19_3/n127 , \add_x_19_3/n126 , \add_x_19_3/n125 ,
         \add_x_19_3/n124 , \add_x_19_3/n123 , \add_x_19_3/n122 ,
         \add_x_19_3/n121 , \add_x_19_3/n120 , \add_x_19_3/n118 ,
         \add_x_19_3/n116 , \add_x_19_3/n113 , \add_x_19_3/n111 ,
         \add_x_19_3/n110 , \add_x_19_3/n106 , \add_x_19_3/n105 ,
         \add_x_19_3/n104 , \add_x_19_3/n103 , \add_x_19_3/n102 ,
         \add_x_19_3/n101 , \add_x_19_3/n100 , \add_x_19_3/n99 ,
         \add_x_19_3/n98 , \add_x_19_3/n97 , \add_x_19_3/n96 ,
         \add_x_19_3/n95 , \add_x_19_3/n94 , \add_x_19_3/n93 ,
         \add_x_19_3/n92 , \add_x_19_3/n91 , \add_x_19_3/n90 ,
         \add_x_19_3/n89 , \add_x_19_3/n88 , \add_x_19_3/n87 ,
         \add_x_19_3/n86 , \add_x_19_3/n85 , \add_x_19_3/n84 ,
         \add_x_19_3/n83 , \add_x_19_3/n82 , \add_x_19_3/n81 ,
         \add_x_19_3/n79 , \add_x_19_3/n78 , \add_x_19_3/n77 ,
         \add_x_19_3/n76 , \add_x_19_3/n75 , \add_x_19_3/n74 ,
         \add_x_19_3/n73 , \add_x_19_3/n72 , \add_x_19_3/n71 ,
         \add_x_19_3/n70 , \add_x_19_3/n69 , \add_x_19_3/n68 ,
         \add_x_19_3/n67 , \add_x_19_3/n66 , \add_x_19_3/n65 ,
         \add_x_19_3/n64 , \add_x_19_3/n63 , \add_x_19_3/n62 ,
         \add_x_19_3/n61 , \add_x_19_3/n60 , \add_x_19_3/n59 ,
         \add_x_19_3/n58 , \add_x_19_3/n56 , \add_x_19_3/n55 ,
         \add_x_19_3/n54 , \add_x_19_3/n53 , \add_x_19_3/n52 ,
         \add_x_19_3/n51 , \add_x_19_3/n50 , \add_x_19_3/n49 ,
         \add_x_19_3/n48 , \add_x_19_3/n47 , \add_x_19_3/n46 ,
         \add_x_19_3/n43 , \add_x_19_3/n42 , \add_x_19_3/n38 ,
         \add_x_19_3/n37 , \add_x_19_3/n36 , \add_x_19_3/n35 ,
         \add_x_19_3/n34 , \add_x_19_3/n30 , \add_x_19_3/n28 ,
         \add_x_19_3/n27 , \add_x_19_3/n26 , \add_x_19_3/n24 ,
         \add_x_19_3/n22 , \add_x_19_3/n18 , \add_x_19_3/n17 ,
         \add_x_19_3/n13 , \add_x_19_3/n11 , \add_x_19_3/n7 , \add_x_19_3/n4 ,
         \add_x_19_5/n222 , \add_x_19_5/n220 , \add_x_19_5/n219 ,
         \add_x_19_5/n214 , \add_x_19_5/n213 , \add_x_19_5/n210 ,
         \add_x_19_5/n207 , \add_x_19_5/n206 , \add_x_19_5/n202 ,
         \add_x_19_5/n198 , \add_x_19_5/n195 , \add_x_19_5/n191 ,
         \add_x_19_5/n189 , \add_x_19_5/n188 , \add_x_19_5/n187 ,
         \add_x_19_5/n186 , \add_x_19_5/n185 , \add_x_19_5/n184 ,
         \add_x_19_5/n183 , \add_x_19_5/n182 , \add_x_19_5/n181 ,
         \add_x_19_5/n180 , \add_x_19_5/n179 , \add_x_19_5/n178 ,
         \add_x_19_5/n176 , \add_x_19_5/n175 , \add_x_19_5/n171 ,
         \add_x_19_5/n170 , \add_x_19_5/n169 , \add_x_19_5/n168 ,
         \add_x_19_5/n167 , \add_x_19_5/n166 , \add_x_19_5/n165 ,
         \add_x_19_5/n163 , \add_x_19_5/n162 , \add_x_19_5/n161 ,
         \add_x_19_5/n160 , \add_x_19_5/n159 , \add_x_19_5/n158 ,
         \add_x_19_5/n157 , \add_x_19_5/n156 , \add_x_19_5/n155 ,
         \add_x_19_5/n154 , \add_x_19_5/n153 , \add_x_19_5/n152 ,
         \add_x_19_5/n151 , \add_x_19_5/n150 , \add_x_19_5/n149 ,
         \add_x_19_5/n148 , \add_x_19_5/n147 , \add_x_19_5/n146 ,
         \add_x_19_5/n145 , \add_x_19_5/n144 , \add_x_19_5/n140 ,
         \add_x_19_5/n139 , \add_x_19_5/n138 , \add_x_19_5/n137 ,
         \add_x_19_5/n136 , \add_x_19_5/n135 , \add_x_19_5/n134 ,
         \add_x_19_5/n133 , \add_x_19_5/n132 , \add_x_19_5/n131 ,
         \add_x_19_5/n130 , \add_x_19_5/n129 , \add_x_19_5/n128 ,
         \add_x_19_5/n127 , \add_x_19_5/n126 , \add_x_19_5/n125 ,
         \add_x_19_5/n124 , \add_x_19_5/n123 , \add_x_19_5/n121 ,
         \add_x_19_5/n120 , \add_x_19_5/n118 , \add_x_19_5/n116 ,
         \add_x_19_5/n113 , \add_x_19_5/n112 , \add_x_19_5/n111 ,
         \add_x_19_5/n110 , \add_x_19_5/n109 , \add_x_19_5/n107 ,
         \add_x_19_5/n106 , \add_x_19_5/n105 , \add_x_19_5/n104 ,
         \add_x_19_5/n103 , \add_x_19_5/n102 , \add_x_19_5/n101 ,
         \add_x_19_5/n100 , \add_x_19_5/n98 , \add_x_19_5/n97 ,
         \add_x_19_5/n96 , \add_x_19_5/n95 , \add_x_19_5/n94 ,
         \add_x_19_5/n93 , \add_x_19_5/n92 , \add_x_19_5/n91 ,
         \add_x_19_5/n90 , \add_x_19_5/n89 , \add_x_19_5/n88 ,
         \add_x_19_5/n87 , \add_x_19_5/n86 , \add_x_19_5/n85 ,
         \add_x_19_5/n84 , \add_x_19_5/n83 , \add_x_19_5/n82 ,
         \add_x_19_5/n81 , \add_x_19_5/n79 , \add_x_19_5/n78 ,
         \add_x_19_5/n76 , \add_x_19_5/n74 , \add_x_19_5/n73 ,
         \add_x_19_5/n72 , \add_x_19_5/n71 , \add_x_19_5/n70 ,
         \add_x_19_5/n69 , \add_x_19_5/n68 , \add_x_19_5/n67 ,
         \add_x_19_5/n66 , \add_x_19_5/n65 , \add_x_19_5/n64 ,
         \add_x_19_5/n63 , \add_x_19_5/n62 , \add_x_19_5/n61 ,
         \add_x_19_5/n60 , \add_x_19_5/n59 , \add_x_19_5/n58 ,
         \add_x_19_5/n56 , \add_x_19_5/n55 , \add_x_19_5/n53 ,
         \add_x_19_5/n52 , \add_x_19_5/n51 , \add_x_19_5/n50 ,
         \add_x_19_5/n49 , \add_x_19_5/n48 , \add_x_19_5/n46 ,
         \add_x_19_5/n43 , \add_x_19_5/n42 , \add_x_19_5/n37 ,
         \add_x_19_5/n36 , \add_x_19_5/n31 , \add_x_19_5/n29 ,
         \add_x_19_5/n28 , \add_x_19_5/n23 , \add_x_19_5/n22 ,
         \add_x_19_5/n19 , \add_x_19_5/n16 , \add_x_19_5/n15 ,
         \add_x_19_5/n11 , \add_x_19_5/n7 , \add_x_19_5/n4 , \add_x_19_0/n219 ,
         \add_x_19_0/n215 , \add_x_19_0/n213 , \add_x_19_0/n210 ,
         \add_x_19_0/n208 , \add_x_19_0/n207 , \add_x_19_0/n206 ,
         \add_x_19_0/n204 , \add_x_19_0/n202 , \add_x_19_0/n198 ,
         \add_x_19_0/n195 , \add_x_19_0/n191 , \add_x_19_0/n189 ,
         \add_x_19_0/n188 , \add_x_19_0/n187 , \add_x_19_0/n186 ,
         \add_x_19_0/n185 , \add_x_19_0/n184 , \add_x_19_0/n182 ,
         \add_x_19_0/n181 , \add_x_19_0/n178 , \add_x_19_0/n177 ,
         \add_x_19_0/n176 , \add_x_19_0/n175 , \add_x_19_0/n171 ,
         \add_x_19_0/n170 , \add_x_19_0/n169 , \add_x_19_0/n168 ,
         \add_x_19_0/n167 , \add_x_19_0/n166 , \add_x_19_0/n165 ,
         \add_x_19_0/n163 , \add_x_19_0/n162 , \add_x_19_0/n156 ,
         \add_x_19_0/n155 , \add_x_19_0/n154 , \add_x_19_0/n152 ,
         \add_x_19_0/n151 , \add_x_19_0/n150 , \add_x_19_0/n149 ,
         \add_x_19_0/n148 , \add_x_19_0/n147 , \add_x_19_0/n146 ,
         \add_x_19_0/n145 , \add_x_19_0/n144 , \add_x_19_0/n140 ,
         \add_x_19_0/n139 , \add_x_19_0/n138 , \add_x_19_0/n137 ,
         \add_x_19_0/n136 , \add_x_19_0/n135 , \add_x_19_0/n134 ,
         \add_x_19_0/n133 , \add_x_19_0/n132 , \add_x_19_0/n131 ,
         \add_x_19_0/n130 , \add_x_19_0/n129 , \add_x_19_0/n128 ,
         \add_x_19_0/n127 , \add_x_19_0/n126 , \add_x_19_0/n125 ,
         \add_x_19_0/n124 , \add_x_19_0/n123 , \add_x_19_0/n122 ,
         \add_x_19_0/n121 , \add_x_19_0/n120 , \add_x_19_0/n118 ,
         \add_x_19_0/n112 , \add_x_19_0/n111 , \add_x_19_0/n110 ,
         \add_x_19_0/n109 , \add_x_19_0/n107 , \add_x_19_0/n106 ,
         \add_x_19_0/n105 , \add_x_19_0/n104 , \add_x_19_0/n103 ,
         \add_x_19_0/n102 , \add_x_19_0/n101 , \add_x_19_0/n100 ,
         \add_x_19_0/n99 , \add_x_19_0/n98 , \add_x_19_0/n97 ,
         \add_x_19_0/n96 , \add_x_19_0/n95 , \add_x_19_0/n94 ,
         \add_x_19_0/n93 , \add_x_19_0/n91 , \add_x_19_0/n90 ,
         \add_x_19_0/n89 , \add_x_19_0/n88 , \add_x_19_0/n87 ,
         \add_x_19_0/n86 , \add_x_19_0/n85 , \add_x_19_0/n84 ,
         \add_x_19_0/n82 , \add_x_19_0/n81 , \add_x_19_0/n79 ,
         \add_x_19_0/n78 , \add_x_19_0/n76 , \add_x_19_0/n74 ,
         \add_x_19_0/n73 , \add_x_19_0/n72 , \add_x_19_0/n69 ,
         \add_x_19_0/n68 , \add_x_19_0/n67 , \add_x_19_0/n66 ,
         \add_x_19_0/n65 , \add_x_19_0/n64 , \add_x_19_0/n63 ,
         \add_x_19_0/n62 , \add_x_19_0/n61 , \add_x_19_0/n60 ,
         \add_x_19_0/n59 , \add_x_19_0/n58 , \add_x_19_0/n56 ,
         \add_x_19_0/n55 , \add_x_19_0/n54 , \add_x_19_0/n53 ,
         \add_x_19_0/n52 , \add_x_19_0/n51 , \add_x_19_0/n50 ,
         \add_x_19_0/n49 , \add_x_19_0/n48 , \add_x_19_0/n47 ,
         \add_x_19_0/n46 , \add_x_19_0/n45 , \add_x_19_0/n44 ,
         \add_x_19_0/n43 , \add_x_19_0/n42 , \add_x_19_0/n38 ,
         \add_x_19_0/n37 , \add_x_19_0/n36 , \add_x_19_0/n35 ,
         \add_x_19_0/n34 , \add_x_19_0/n28 , \add_x_19_0/n24 ,
         \add_x_19_0/n22 , \add_x_19_0/n19 , \add_x_19_0/n17 ,
         \add_x_19_0/n15 , \add_x_19_0/n13 , \add_x_19_0/n11 , \add_x_19_0/n7 ,
         \add_x_19_0/n4 , \add_x_19_0/n1 , \DP_OP_159_297_3515/n1138 ,
         \DP_OP_159_297_3515/n1133 , \DP_OP_159_297_3515/n1128 ,
         \DP_OP_159_297_3515/n1074 , \DP_OP_159_297_3515/n1069 ,
         \DP_OP_159_297_3515/n1064 , \DP_OP_159_297_3515/n1063 ,
         \DP_OP_159_297_3515/n1057 , \DP_OP_159_297_3515/n1052 ,
         \DP_OP_159_297_3515/n1051 , \DP_OP_159_297_3515/n1044 ,
         \DP_OP_159_297_3515/n1039 , \DP_OP_159_297_3515/n1031 ,
         \DP_OP_159_297_3515/n1026 , \DP_OP_159_297_3515/n1025 ,
         \DP_OP_159_297_3515/n1024 , \DP_OP_159_297_3515/n1018 ,
         \DP_OP_159_297_3515/n1017 , \DP_OP_159_297_3515/n1012 ,
         \DP_OP_159_297_3515/n1011 , \DP_OP_159_297_3515/n1010 ,
         \DP_OP_159_297_3515/n1004 , \DP_OP_159_297_3515/n1003 ,
         \DP_OP_159_297_3515/n999 , \DP_OP_159_297_3515/n998 ,
         \DP_OP_159_297_3515/n997 , \DP_OP_159_297_3515/n996 ,
         \DP_OP_159_297_3515/n991 , \DP_OP_159_297_3515/n990 ,
         \DP_OP_159_297_3515/n989 , \DP_OP_159_297_3515/n976 ,
         \DP_OP_159_297_3515/n971 , \DP_OP_159_297_3515/n964 ,
         \DP_OP_159_297_3515/n963 , \DP_OP_159_297_3515/n959 ,
         \DP_OP_159_297_3515/n957 , \DP_OP_159_297_3515/n956 ,
         \DP_OP_159_297_3515/n955 , \DP_OP_159_297_3515/n950 ,
         \DP_OP_159_297_3515/n949 , \DP_OP_159_297_3515/n948 ,
         \DP_OP_159_297_3515/n944 , \DP_OP_159_297_3515/n943 ,
         \DP_OP_159_297_3515/n936 , \DP_OP_159_297_3515/n935 ,
         \DP_OP_159_297_3515/n934 , \DP_OP_159_297_3515/n931 ,
         \DP_OP_159_297_3515/n930 , \DP_OP_159_297_3515/n928 ,
         \DP_OP_159_297_3515/n927 , \DP_OP_159_297_3515/n921 ,
         \DP_OP_159_297_3515/n920 , \DP_OP_159_297_3515/n916 ,
         \DP_OP_159_297_3515/n915 , \DP_OP_159_297_3515/n914 ,
         \DP_OP_159_297_3515/n913 , \DP_OP_159_297_3515/n908 ,
         \DP_OP_159_297_3515/n907 , \DP_OP_159_297_3515/n906 ,
         \DP_OP_159_297_3515/n902 , \DP_OP_159_297_3515/n894 ,
         \DP_OP_159_297_3515/n893 , \DP_OP_159_297_3515/n892 ,
         \DP_OP_159_297_3515/n887 , \DP_OP_159_297_3515/n886 ,
         \DP_OP_159_297_3515/n885 , \DP_OP_159_297_3515/n880 ,
         \DP_OP_159_297_3515/n879 , \DP_OP_159_297_3515/n878 ,
         \DP_OP_159_297_3515/n877 , \DP_OP_159_297_3515/n876 ,
         \DP_OP_159_297_3515/n875 , \DP_OP_159_297_3515/n873 ,
         \DP_OP_159_297_3515/n871 , \DP_OP_159_297_3515/n870 ,
         \DP_OP_159_297_3515/n869 , \DP_OP_159_297_3515/n868 ,
         \DP_OP_159_297_3515/n867 , \DP_OP_159_297_3515/n862 ,
         \DP_OP_159_297_3515/n852 , \DP_OP_159_297_3515/n815 ,
         \DP_OP_159_297_3515/n778 , \DP_OP_159_297_3515/n776 ,
         \DP_OP_159_297_3515/n774 , \DP_OP_159_297_3515/n768 ,
         \DP_OP_159_297_3515/n766 , \DP_OP_159_297_3515/n764 ,
         \DP_OP_159_297_3515/n758 , \DP_OP_159_297_3515/n742 ,
         \DP_OP_159_297_3515/n740 , \DP_OP_159_297_3515/n737 ,
         \DP_OP_159_297_3515/n730 , \DP_OP_159_297_3515/n728 ,
         \DP_OP_159_297_3515/n726 , \DP_OP_159_297_3515/n723 ,
         \DP_OP_159_297_3515/n714 , \DP_OP_159_297_3515/n712 ,
         \DP_OP_159_297_3515/n705 , \DP_OP_159_297_3515/n694 ,
         \DP_OP_159_297_3515/n692 , \DP_OP_159_297_3515/n690 ,
         \DP_OP_159_297_3515/n688 , \DP_OP_159_297_3515/n685 ,
         \DP_OP_159_297_3515/n674 , \DP_OP_159_297_3515/n672 ,
         \DP_OP_159_297_3515/n650 , \DP_OP_159_297_3515/n648 ,
         \DP_OP_159_297_3515/n646 , \DP_OP_159_297_3515/n638 ,
         \DP_OP_159_297_3515/n625 , \DP_OP_159_297_3515/n623 ,
         \DP_OP_159_297_3515/n610 , \DP_OP_159_297_3515/n593 ,
         \DP_OP_159_297_3515/n591 , \DP_OP_159_297_3515/n589 ,
         \DP_OP_159_297_3515/n587 , \DP_OP_159_297_3515/n160 ,
         \DP_OP_159_297_3515/n1 , \DP_OP_158_296_6262/n2060 ,
         \DP_OP_158_296_6262/n2054 , \DP_OP_158_296_6262/n2051 ,
         \DP_OP_158_296_6262/n2048 , \DP_OP_158_296_6262/n2034 ,
         \DP_OP_158_296_6262/n2020 , \DP_OP_158_296_6262/n2015 ,
         \DP_OP_158_296_6262/n2011 , \DP_OP_158_296_6262/n2010 ,
         \DP_OP_158_296_6262/n2004 , \DP_OP_158_296_6262/n1999 ,
         \DP_OP_158_296_6262/n1998 , \DP_OP_158_296_6262/n1991 ,
         \DP_OP_158_296_6262/n1987 , \DP_OP_158_296_6262/n1978 ,
         \DP_OP_158_296_6262/n1973 , \DP_OP_158_296_6262/n1972 ,
         \DP_OP_158_296_6262/n1971 , \DP_OP_158_296_6262/n1966 ,
         \DP_OP_158_296_6262/n1965 , \DP_OP_158_296_6262/n1964 ,
         \DP_OP_158_296_6262/n1959 , \DP_OP_158_296_6262/n1958 ,
         \DP_OP_158_296_6262/n1957 , \DP_OP_158_296_6262/n1952 ,
         \DP_OP_158_296_6262/n1951 , \DP_OP_158_296_6262/n1950 ,
         \DP_OP_158_296_6262/n1946 , \DP_OP_158_296_6262/n1945 ,
         \DP_OP_158_296_6262/n1944 , \DP_OP_158_296_6262/n1943 ,
         \DP_OP_158_296_6262/n1938 , \DP_OP_158_296_6262/n1937 ,
         \DP_OP_158_296_6262/n1936 , \DP_OP_158_296_6262/n1918 ,
         \DP_OP_158_296_6262/n1917 , \DP_OP_158_296_6262/n1916 ,
         \DP_OP_158_296_6262/n1911 , \DP_OP_158_296_6262/n1910 ,
         \DP_OP_158_296_6262/n1909 , \DP_OP_158_296_6262/n1904 ,
         \DP_OP_158_296_6262/n1903 , \DP_OP_158_296_6262/n1897 ,
         \DP_OP_158_296_6262/n1896 , \DP_OP_158_296_6262/n1895 ,
         \DP_OP_158_296_6262/n1890 , \DP_OP_158_296_6262/n1881 ,
         \DP_OP_158_296_6262/n1877 , \DP_OP_158_296_6262/n1875 ,
         \DP_OP_158_296_6262/n1874 , \DP_OP_158_296_6262/n1869 ,
         \DP_OP_158_296_6262/n1863 , \DP_OP_158_296_6262/n1862 ,
         \DP_OP_158_296_6262/n1855 , \DP_OP_158_296_6262/n1854 ,
         \DP_OP_158_296_6262/n1849 , \DP_OP_158_296_6262/n1848 ,
         \DP_OP_158_296_6262/n1847 , \DP_OP_158_296_6262/n1837 ,
         \DP_OP_158_296_6262/n1834 , \DP_OP_158_296_6262/n1833 ,
         \DP_OP_158_296_6262/n1830 , \DP_OP_158_296_6262/n1829 ,
         \DP_OP_158_296_6262/n1828 , \DP_OP_158_296_6262/n1827 ,
         \DP_OP_158_296_6262/n1826 , \DP_OP_158_296_6262/n1792 ,
         \DP_OP_158_296_6262/n1791 , \DP_OP_158_296_6262/n855 ,
         \DP_OP_158_296_6262/n841 , \DP_OP_158_296_6262/n838 ,
         \DP_OP_158_296_6262/n833 , \DP_OP_158_296_6262/n829 ,
         \DP_OP_158_296_6262/n375 , \DP_OP_158_296_6262/n373 ,
         \DP_OP_158_296_6262/n371 , \DP_OP_158_296_6262/n365 ,
         \DP_OP_158_296_6262/n349 , \DP_OP_158_296_6262/n347 ,
         \DP_OP_158_296_6262/n329 , \DP_OP_158_296_6262/n322 ,
         \DP_OP_158_296_6262/n320 , \DP_OP_158_296_6262/n318 ,
         \DP_OP_158_296_6262/n315 , \DP_OP_158_296_6262/n306 ,
         \DP_OP_158_296_6262/n304 , \DP_OP_158_296_6262/n297 ,
         \DP_OP_158_296_6262/n286 , \DP_OP_158_296_6262/n284 ,
         \DP_OP_158_296_6262/n282 , \DP_OP_158_296_6262/n280 ,
         \DP_OP_158_296_6262/n277 , \DP_OP_158_296_6262/n266 ,
         \DP_OP_158_296_6262/n264 , \DP_OP_158_296_6262/n255 ,
         \DP_OP_158_296_6262/n242 , \DP_OP_158_296_6262/n240 ,
         \DP_OP_158_296_6262/n238 , \DP_OP_158_296_6262/n230 ,
         \DP_OP_158_296_6262/n217 , \DP_OP_158_296_6262/n215 ,
         \DP_OP_158_296_6262/n202 , \DP_OP_158_296_6262/n185 ,
         \DP_OP_158_296_6262/n183 , \DP_OP_158_296_6262/n181 ,
         \DP_OP_158_296_6262/n179 , \DP_OP_158_296_6262/n174 ,
         \DP_OP_158_296_6262/n161 , \DP_OP_158_296_6262/n159 ,
         \DP_OP_158_296_6262/n148 , \DP_OP_158_296_6262/n133 ,
         \DP_OP_158_296_6262/n131 , \DP_OP_158_296_6262/n129 ,
         \DP_OP_158_296_6262/n119 , \DP_OP_158_296_6262/n104 ,
         \DP_OP_158_296_6262/n102 , \DP_OP_158_296_6262/n87 ,
         \DP_OP_158_296_6262/n68 , \DP_OP_158_296_6262/n66 ,
         \DP_OP_158_296_6262/n64 , \DP_OP_158_296_6262/n62 ,
         \DP_OP_158_296_6262/n54 , \DP_OP_158_296_6262/n39 ,
         \DP_OP_158_296_6262/n37 , \DP_OP_158_296_6262/n18 ,
         \DP_OP_158_296_6262/n5 , \DP_OP_158_296_6262/n3 , \add_x_22_4/n121 ,
         \add_x_22_4/n119 , \add_x_22_4/n118 , \add_x_22_4/n117 ,
         \add_x_22_4/n115 , \add_x_22_4/n112 , \add_x_22_4/n111 ,
         \add_x_22_4/n110 , \add_x_22_4/n109 , \add_x_22_4/n106 ,
         \add_x_22_4/n105 , \add_x_22_4/n103 , \add_x_22_4/n102 ,
         \add_x_22_4/n101 , \add_x_22_4/n99 , \add_x_22_4/n98 ,
         \add_x_22_4/n94 , \add_x_22_4/n93 , \add_x_22_4/n92 ,
         \add_x_22_4/n90 , \add_x_22_4/n87 , \add_x_22_4/n85 ,
         \add_x_22_4/n84 , \add_x_22_4/n81 , \add_x_22_4/n80 ,
         \add_x_22_4/n78 , \add_x_22_4/n77 , \add_x_22_4/n76 ,
         \add_x_22_4/n75 , \add_x_22_4/n74 , \add_x_22_4/n71 ,
         \add_x_22_4/n69 , \add_x_22_4/n68 , \add_x_22_4/n67 ,
         \add_x_22_4/n65 , \add_x_22_4/n64 , \add_x_22_4/n59 ,
         \add_x_22_4/n58 , \add_x_22_4/n57 , \add_x_22_4/n54 ,
         \add_x_22_4/n51 , \add_x_22_4/n50 , \add_x_22_4/n47 ,
         \add_x_22_4/n46 , \add_x_22_4/n44 , \add_x_22_4/n43 ,
         \add_x_22_4/n42 , \add_x_22_4/n41 , \add_x_22_4/n35 ,
         \add_x_22_4/n34 , \add_x_22_4/n33 , \add_x_22_4/n30 ,
         \add_x_22_4/n28 , \add_x_22_4/n27 , \add_x_22_4/n26 ,
         \add_x_22_4/n24 , \add_x_22_4/n23 , \add_x_22_4/n20 ,
         \add_x_22_4/n17 , \add_x_22_4/n16 , \add_x_22_4/n15 ,
         \add_x_22_4/n10 , \add_x_22_4/n9 , \add_x_22_4/n8 , \add_x_22_4/n7 ,
         \add_x_22_4/n2 , \add_x_22_4/n1 , \add_x_22_1/n121 ,
         \add_x_22_1/n119 , \add_x_22_1/n118 , \add_x_22_1/n117 ,
         \add_x_22_1/n115 , \add_x_22_1/n114 , \add_x_22_1/n112 ,
         \add_x_22_1/n111 , \add_x_22_1/n110 , \add_x_22_1/n109 ,
         \add_x_22_1/n103 , \add_x_22_1/n102 , \add_x_22_1/n99 ,
         \add_x_22_1/n98 , \add_x_22_1/n96 , \add_x_22_1/n95 ,
         \add_x_22_1/n94 , \add_x_22_1/n93 , \add_x_22_1/n92 ,
         \add_x_22_1/n90 , \add_x_22_1/n89 , \add_x_22_1/n87 ,
         \add_x_22_1/n85 , \add_x_22_1/n84 , \add_x_22_1/n78 ,
         \add_x_22_1/n77 , \add_x_22_1/n76 , \add_x_22_1/n75 ,
         \add_x_22_1/n74 , \add_x_22_1/n72 , \add_x_22_1/n71 ,
         \add_x_22_1/n69 , \add_x_22_1/n68 , \add_x_22_1/n67 ,
         \add_x_22_1/n65 , \add_x_22_1/n64 , \add_x_22_1/n59 ,
         \add_x_22_1/n58 , \add_x_22_1/n57 , \add_x_22_1/n54 ,
         \add_x_22_1/n53 , \add_x_22_1/n51 , \add_x_22_1/n50 ,
         \add_x_22_1/n47 , \add_x_22_1/n44 , \add_x_22_1/n43 ,
         \add_x_22_1/n42 , \add_x_22_1/n41 , \add_x_22_1/n38 ,
         \add_x_22_1/n35 , \add_x_22_1/n34 , \add_x_22_1/n31 ,
         \add_x_22_1/n30 , \add_x_22_1/n28 , \add_x_22_1/n27 ,
         \add_x_22_1/n26 , \add_x_22_1/n24 , \add_x_22_1/n23 ,
         \add_x_22_1/n20 , \add_x_22_1/n17 , \add_x_22_1/n16 ,
         \add_x_22_1/n15 , \add_x_22_1/n10 , \add_x_22_1/n9 , \add_x_22_1/n8 ,
         \add_x_22_1/n7 , \add_x_22_1/n5 , \add_x_22_1/n4 , \add_x_22_1/n3 ,
         \add_x_22_1/n2 , \add_x_22_1/n1 , \add_x_22_5/n121 ,
         \add_x_22_5/n119 , \add_x_22_5/n118 , \add_x_22_5/n117 ,
         \add_x_22_5/n115 , \add_x_22_5/n114 , \add_x_22_5/n112 ,
         \add_x_22_5/n111 , \add_x_22_5/n110 , \add_x_22_5/n109 ,
         \add_x_22_5/n106 , \add_x_22_5/n103 , \add_x_22_5/n102 ,
         \add_x_22_5/n101 , \add_x_22_5/n99 , \add_x_22_5/n94 ,
         \add_x_22_5/n93 , \add_x_22_5/n92 , \add_x_22_5/n90 ,
         \add_x_22_5/n89 , \add_x_22_5/n87 , \add_x_22_5/n85 ,
         \add_x_22_5/n84 , \add_x_22_5/n81 , \add_x_22_5/n80 ,
         \add_x_22_5/n78 , \add_x_22_5/n77 , \add_x_22_5/n76 ,
         \add_x_22_5/n75 , \add_x_22_5/n74 , \add_x_22_5/n72 ,
         \add_x_22_5/n71 , \add_x_22_5/n69 , \add_x_22_5/n68 ,
         \add_x_22_5/n67 , \add_x_22_5/n64 , \add_x_22_5/n59 ,
         \add_x_22_5/n58 , \add_x_22_5/n57 , \add_x_22_5/n54 ,
         \add_x_22_5/n53 , \add_x_22_5/n51 , \add_x_22_5/n50 ,
         \add_x_22_5/n49 , \add_x_22_5/n47 , \add_x_22_5/n44 ,
         \add_x_22_5/n43 , \add_x_22_5/n42 , \add_x_22_5/n41 ,
         \add_x_22_5/n35 , \add_x_22_5/n34 , \add_x_22_5/n33 ,
         \add_x_22_5/n31 , \add_x_22_5/n26 , \add_x_22_5/n24 ,
         \add_x_22_5/n23 , \add_x_22_5/n20 , \add_x_22_5/n17 ,
         \add_x_22_5/n16 , \add_x_22_5/n15 , \add_x_22_5/n13 ,
         \add_x_22_5/n10 , \add_x_22_5/n9 , \add_x_22_5/n8 , \add_x_22_5/n5 ,
         \add_x_22_5/n4 , \add_x_22_5/n3 , \add_x_22_5/n2 , \add_x_22_5/n1 ,
         \add_x_22_3/n119 , \add_x_22_3/n118 , \add_x_22_3/n115 ,
         \add_x_22_3/n114 , \add_x_22_3/n112 , \add_x_22_3/n111 ,
         \add_x_22_3/n110 , \add_x_22_3/n109 , \add_x_22_3/n106 ,
         \add_x_22_3/n105 , \add_x_22_3/n103 , \add_x_22_3/n102 ,
         \add_x_22_3/n101 , \add_x_22_3/n98 , \add_x_22_3/n94 ,
         \add_x_22_3/n93 , \add_x_22_3/n92 , \add_x_22_3/n90 ,
         \add_x_22_3/n89 , \add_x_22_3/n87 , \add_x_22_3/n85 ,
         \add_x_22_3/n84 , \add_x_22_3/n81 , \add_x_22_3/n80 ,
         \add_x_22_3/n78 , \add_x_22_3/n77 , \add_x_22_3/n76 ,
         \add_x_22_3/n75 , \add_x_22_3/n72 , \add_x_22_3/n71 ,
         \add_x_22_3/n69 , \add_x_22_3/n68 , \add_x_22_3/n59 ,
         \add_x_22_3/n58 , \add_x_22_3/n57 , \add_x_22_3/n54 ,
         \add_x_22_3/n51 , \add_x_22_3/n50 , \add_x_22_3/n47 ,
         \add_x_22_3/n44 , \add_x_22_3/n43 , \add_x_22_3/n42 ,
         \add_x_22_3/n41 , \add_x_22_3/n35 , \add_x_22_3/n34 ,
         \add_x_22_3/n31 , \add_x_22_3/n30 , \add_x_22_3/n28 ,
         \add_x_22_3/n27 , \add_x_22_3/n26 , \add_x_22_3/n24 ,
         \add_x_22_3/n23 , \add_x_22_3/n22 , \add_x_22_3/n20 ,
         \add_x_22_3/n19 , \add_x_22_3/n17 , \add_x_22_3/n16 ,
         \add_x_22_3/n15 , \add_x_22_3/n13 , \add_x_22_3/n10 , \add_x_22_3/n9 ,
         \add_x_22_3/n8 , \add_x_22_3/n7 , \add_x_22_3/n2 , \add_x_22_3/n1 ,
         \add_x_22_2/n121 , \add_x_22_2/n119 , \add_x_22_2/n118 ,
         \add_x_22_2/n117 , \add_x_22_2/n114 , \add_x_22_2/n112 ,
         \add_x_22_2/n111 , \add_x_22_2/n110 , \add_x_22_2/n109 ,
         \add_x_22_2/n106 , \add_x_22_2/n105 , \add_x_22_2/n103 ,
         \add_x_22_2/n102 , \add_x_22_2/n101 , \add_x_22_2/n99 ,
         \add_x_22_2/n98 , \add_x_22_2/n94 , \add_x_22_2/n93 ,
         \add_x_22_2/n92 , \add_x_22_2/n90 , \add_x_22_2/n87 ,
         \add_x_22_2/n85 , \add_x_22_2/n81 , \add_x_22_2/n80 ,
         \add_x_22_2/n78 , \add_x_22_2/n77 , \add_x_22_2/n76 ,
         \add_x_22_2/n75 , \add_x_22_2/n74 , \add_x_22_2/n72 ,
         \add_x_22_2/n71 , \add_x_22_2/n69 , \add_x_22_2/n68 ,
         \add_x_22_2/n64 , \add_x_22_2/n59 , \add_x_22_2/n58 ,
         \add_x_22_2/n54 , \add_x_22_2/n53 , \add_x_22_2/n51 ,
         \add_x_22_2/n50 , \add_x_22_2/n47 , \add_x_22_2/n46 ,
         \add_x_22_2/n44 , \add_x_22_2/n43 , \add_x_22_2/n42 ,
         \add_x_22_2/n41 , \add_x_22_2/n38 , \add_x_22_2/n35 ,
         \add_x_22_2/n34 , \add_x_22_2/n31 , \add_x_22_2/n30 ,
         \add_x_22_2/n26 , \add_x_22_2/n24 , \add_x_22_2/n23 ,
         \add_x_22_2/n17 , \add_x_22_2/n16 , \add_x_22_2/n15 ,
         \add_x_22_2/n12 , \add_x_22_2/n10 , \add_x_22_2/n9 , \add_x_22_2/n8 ,
         \add_x_22_2/n2 , \add_x_22_2/n1 , \add_x_22_0/n121 ,
         \add_x_22_0/n119 , \add_x_22_0/n118 , \add_x_22_0/n117 ,
         \add_x_22_0/n115 , \add_x_22_0/n114 , \add_x_22_0/n112 ,
         \add_x_22_0/n111 , \add_x_22_0/n110 , \add_x_22_0/n109 ,
         \add_x_22_0/n106 , \add_x_22_0/n105 , \add_x_22_0/n103 ,
         \add_x_22_0/n102 , \add_x_22_0/n101 , \add_x_22_0/n99 ,
         \add_x_22_0/n96 , \add_x_22_0/n95 , \add_x_22_0/n94 ,
         \add_x_22_0/n93 , \add_x_22_0/n92 , \add_x_22_0/n90 ,
         \add_x_22_0/n89 , \add_x_22_0/n87 , \add_x_22_0/n85 ,
         \add_x_22_0/n84 , \add_x_22_0/n80 , \add_x_22_0/n78 ,
         \add_x_22_0/n77 , \add_x_22_0/n76 , \add_x_22_0/n75 ,
         \add_x_22_0/n72 , \add_x_22_0/n69 , \add_x_22_0/n68 ,
         \add_x_22_0/n65 , \add_x_22_0/n59 , \add_x_22_0/n58 ,
         \add_x_22_0/n57 , \add_x_22_0/n51 , \add_x_22_0/n50 ,
         \add_x_22_0/n49 , \add_x_22_0/n47 , \add_x_22_0/n44 ,
         \add_x_22_0/n43 , \add_x_22_0/n42 , \add_x_22_0/n41 ,
         \add_x_22_0/n40 , \add_x_22_0/n35 , \add_x_22_0/n34 ,
         \add_x_22_0/n31 , \add_x_22_0/n26 , \add_x_22_0/n24 ,
         \add_x_22_0/n23 , \add_x_22_0/n20 , \add_x_22_0/n17 ,
         \add_x_22_0/n16 , \add_x_22_0/n15 , \add_x_22_0/n13 ,
         \add_x_22_0/n10 , \add_x_22_0/n9 , \add_x_22_0/n8 , \add_x_22_0/n7 ,
         \add_x_22_0/n5 , \add_x_22_0/n4 , \add_x_22_0/n3 , \add_x_22_0/n2 ,
         \add_x_22_0/n1 , \DP_OP_159_297_3515/n1075 ,
         \DP_OP_159_297_3515/n1066 , \DP_OP_158_296_6262/n2056 ,
         \DP_OP_158_296_6262/n1861 , \DP_OP_158_296_6262/n1860 ,
         \add_x_19_4/n50 , \add_x_19_4/n4 , \add_x_19_4/n195 , \add_x_19_4/n7 ,
         \add_x_19_4/n65 , \add_x_19_4/n198 , \add_x_19_4/n71 ,
         \add_x_19_4/n70 , \add_x_19_4/n119 , \add_x_19_4/n117 ,
         \add_x_19_4/n115 , \add_x_19_4/n114 , \add_x_19_4/n40 ,
         \add_x_19_4/n47 , \add_x_19_4/n45 , \add_x_19_4/n44 ,
         \add_x_19_4/n208 , \add_x_19_4/n17 , \add_x_19_4/n122 ,
         \addr_calc/fft_write_calc/counter/N48 , \add_x_22_1/n106 ,
         \DP_OP_159_297_3515/n87 , \DP_OP_159_297_3515/n85 ,
         \DP_OP_159_297_3515/n792 , \DP_OP_159_297_3515/n70 ,
         \DP_OP_159_297_3515/n51 , \DP_OP_159_297_3515/n5 ,
         \DP_OP_159_297_3515/n49 , \DP_OP_159_297_3515/n47 ,
         \DP_OP_159_297_3515/n45 , \DP_OP_159_297_3515/n3 ,
         \DP_OP_159_297_3515/n18 , \DP_OP_159_297_3515/n157 ,
         \DP_OP_159_297_3515/n144 , \DP_OP_159_297_3515/n142 ,
         \DP_OP_159_297_3515/n131 , \DP_OP_159_297_3515/n116 ,
         \DP_OP_159_297_3515/n114 , \DP_OP_159_297_3515/n112 ,
         \DP_OP_159_297_3515/n102 , \DP_OP_159_297_3515/n942 ,
         \DP_OP_159_297_3515/n941 , \DP_OP_159_297_3515/n861 ,
         \DP_OP_158_296_6262/n1891 , \DP_OP_158_296_6262/n1883 ,
         \DP_OP_158_296_6262/n1882 , \DP_OP_158_296_6262/n1906 ,
         \DP_OP_158_296_6262/n1878 , \add_x_19_0/n119 , \add_x_19_0/n117 ,
         \add_x_19_0/n115 , \add_x_19_0/n114 , \add_x_19_0/n161 ,
         \add_x_19_0/n159 , \add_x_19_0/n158 , \DP_OP_158_296_6262/n998 ,
         \DP_OP_158_296_6262/n996 , \DP_OP_158_296_6262/n981 ,
         \DP_OP_158_296_6262/n962 , \DP_OP_158_296_6262/n960 ,
         \DP_OP_158_296_6262/n958 , \DP_OP_158_296_6262/n956 ,
         \DP_OP_158_296_6262/n948 , \DP_OP_158_296_6262/n933 ,
         \DP_OP_158_296_6262/n931 , \DP_OP_158_296_6262/n912 ,
         \DP_OP_158_296_6262/n899 , \DP_OP_158_296_6262/n897 ,
         \DP_OP_158_296_6262/n895 , \DP_OP_158_296_6262/n1269 ,
         \DP_OP_158_296_6262/n1267 , \DP_OP_158_296_6262/n1265 ,
         \DP_OP_158_296_6262/n1259 , \DP_OP_158_296_6262/n1243 ,
         \DP_OP_158_296_6262/n1241 , \DP_OP_158_296_6262/n1223 ,
         \DP_OP_158_296_6262/n1216 , \DP_OP_158_296_6262/n1214 ,
         \DP_OP_158_296_6262/n1212 , \DP_OP_158_296_6262/n1209 ,
         \DP_OP_158_296_6262/n1200 , \DP_OP_158_296_6262/n1198 ,
         \DP_OP_158_296_6262/n1191 , \DP_OP_158_296_6262/n1180 ,
         \DP_OP_158_296_6262/n1178 , \DP_OP_158_296_6262/n1176 ,
         \DP_OP_158_296_6262/n1174 , \DP_OP_158_296_6262/n1171 ,
         \DP_OP_158_296_6262/n1160 , \DP_OP_158_296_6262/n1158 ,
         \DP_OP_158_296_6262/n1149 , \DP_OP_158_296_6262/n1136 ,
         \DP_OP_158_296_6262/n1134 , \DP_OP_158_296_6262/n1132 ,
         \DP_OP_158_296_6262/n1124 , \DP_OP_158_296_6262/n1111 ,
         \DP_OP_158_296_6262/n1109 , \DP_OP_158_296_6262/n1079 ,
         \DP_OP_158_296_6262/n1077 , \DP_OP_158_296_6262/n1075 ,
         \DP_OP_158_296_6262/n1073 , \DP_OP_158_296_6262/n1071 ,
         \DP_OP_158_296_6262/n1068 , \DP_OP_158_296_6262/n1055 ,
         \DP_OP_158_296_6262/n1053 , \DP_OP_158_296_6262/n1042 ,
         \DP_OP_158_296_6262/n1027 , \DP_OP_158_296_6262/n1025 ,
         \DP_OP_158_296_6262/n1023 , \DP_OP_158_296_6262/n1013 ,
         \DP_OP_158_296_6262/n1842 , \DP_OP_158_296_6262/n1841 ,
         \DP_OP_158_296_6262/n1840 , \DP_OP_158_296_6262/n1850 ,
         \add_x_19_3/n9 , \add_x_19_3/n80 , \add_x_19_3/n200 ,
         \add_x_19_5/n35 , \add_x_19_5/n34 , \add_x_19_5/n1 ,
         \add_x_19_4/n161 , \add_x_19_4/n159 , \add_x_19_4/n158 ,
         \add_x_19_5/n9 , \add_x_19_5/n80 , \add_x_19_5/n200 ,
         \add_x_19_4/n80 , \add_x_19_4/n200 , \add_x_19_3/n138 ,
         \add_x_19_4/n83 , \add_x_19_4/n92 , \add_x_19_4/n113 ,
         \addr_calc/iir_write_calc/counter/N64 , \add_x_22_5/n38 ,
         \addr_calc/iir_write_calc/counter/N38 , \DP_OP_159_297_3515/n582 ,
         \DP_OP_159_297_3515/n569 , \DP_OP_159_297_3515/n567 ,
         \DP_OP_159_297_3515/n556 , \DP_OP_159_297_3515/n541 ,
         \DP_OP_159_297_3515/n539 , \DP_OP_159_297_3515/n537 ,
         \DP_OP_159_297_3515/n527 , \DP_OP_159_297_3515/n512 ,
         \DP_OP_159_297_3515/n510 , \DP_OP_159_297_3515/n495 ,
         \DP_OP_159_297_3515/n476 , \DP_OP_159_297_3515/n474 ,
         \DP_OP_159_297_3515/n472 , \DP_OP_159_297_3515/n470 ,
         \DP_OP_159_297_3515/n443 , \DP_OP_159_297_3515/n430 ,
         \DP_OP_159_297_3515/n428 , \DP_OP_159_297_3515/n901 ,
         \DP_OP_159_297_3515/n900 , \DP_OP_159_297_3515/n899 ,
         \DP_OP_159_297_3515/n903 , \add_x_19_3/n161 , \add_x_19_3/n159 ,
         \add_x_19_3/n158 , \add_x_19_0/n80 , \add_x_19_0/n200 ,
         \add_x_19_2/n35 , \add_x_19_2/n34 , \add_x_19_2/n1 , \add_x_19_0/n83 ,
         \add_x_19_0/n92 , \add_x_19_0/n113 , \add_x_19_0/n157 ,
         \add_x_19_5/n99 , \add_x_19_5/n204 , \add_x_19_5/n13 ,
         \add_x_19_1/n57 , \add_x_19_1/n5 , \add_x_19_1/n196 ,
         \add_x_19_1/n71 , \add_x_19_1/n70 , \add_x_19_1/n180 ,
         \add_x_19_1/n179 , \add_x_19_3/n180 , \add_x_19_3/n179 ,
         \add_x_19_1/n170 , \add_x_19_0/n57 , \add_x_19_0/n196 ,
         \add_x_19_0/n71 , \add_x_19_0/n70 , \add_x_19_5/n117 ,
         \add_x_19_5/n115 , \add_x_19_5/n114 , \add_x_19_0/n77 ,
         \add_x_19_0/n75 , \add_x_19_2/n47 , \add_x_19_2/n45 ,
         \add_x_19_2/n44 , \add_x_19_2/n138 , \add_x_19_4/n180 ,
         \add_x_19_4/n179 , \add_x_19_2/n38 , \add_x_19_2/n43 ,
         \add_x_19_2/n113 , \add_x_19_2/n136 , \add_x_19_2/n145 ,
         \add_x_19_2/n157 , \add_x_19_2/n160 , \add_x_19_2/n162 ,
         \add_x_19_2/n77 , \add_x_19_2/n75 , \add_x_19_5/n47 ,
         \add_x_19_5/n45 , \add_x_19_5/n44 , \add_x_19_5/n77 ,
         \add_x_19_5/n75 , \add_x_19_1/n9 , \add_x_19_1/n80 ,
         \add_x_19_1/n200 , \addr_calc/iir_read_calc/counter/N64 ,
         \add_x_22_4/n38 , \addr_calc/iir_read_calc/counter/N38 ,
         \DP_OP_159_297_3515/n353 , \DP_OP_159_297_3515/n351 ,
         \DP_OP_159_297_3515/n349 , \DP_OP_159_297_3515/n343 ,
         \DP_OP_159_297_3515/n341 , \DP_OP_159_297_3515/n339 ,
         \DP_OP_159_297_3515/n333 , \DP_OP_159_297_3515/n317 ,
         \DP_OP_159_297_3515/n315 , \DP_OP_159_297_3515/n312 ,
         \DP_OP_159_297_3515/n305 , \DP_OP_159_297_3515/n303 ,
         \DP_OP_159_297_3515/n301 , \DP_OP_159_297_3515/n298 ,
         \DP_OP_159_297_3515/n289 , \DP_OP_159_297_3515/n287 ,
         \DP_OP_159_297_3515/n280 , \DP_OP_159_297_3515/n269 ,
         \DP_OP_159_297_3515/n267 , \DP_OP_159_297_3515/n265 ,
         \DP_OP_159_297_3515/n263 , \DP_OP_159_297_3515/n260 ,
         \DP_OP_159_297_3515/n249 , \DP_OP_159_297_3515/n247 ,
         \DP_OP_159_297_3515/n238 , \DP_OP_159_297_3515/n225 ,
         \DP_OP_159_297_3515/n223 , \DP_OP_159_297_3515/n221 ,
         \DP_OP_159_297_3515/n213 , \DP_OP_159_297_3515/n200 ,
         \DP_OP_159_297_3515/n198 , \DP_OP_159_297_3515/n185 ,
         \DP_OP_159_297_3515/n168 , \DP_OP_159_297_3515/n166 ,
         \DP_OP_159_297_3515/n164 , \DP_OP_159_297_3515/n162 ,
         \DP_OP_159_297_3515/n970 , \DP_OP_159_297_3515/n969 ,
         \DP_OP_159_297_3515/n986 , \DP_OP_159_297_3515/n985 ,
         \DP_OP_159_297_3515/n1041 , \DP_OP_159_297_3515/n1040 ,
         \addr_calc/fir_write_calc/counter/N44 , \add_x_22_3/n121 ,
         \addr_calc/fir_write_calc/counter/N50 , \add_x_22_3/n99 ,
         \addr_calc/fir_write_calc/counter/N53 , \DP_OP_158_296_6262/n1716 ,
         \DP_OP_158_296_6262/n1714 , \DP_OP_158_296_6262/n1712 ,
         \DP_OP_158_296_6262/n1706 , \DP_OP_158_296_6262/n1690 ,
         \DP_OP_158_296_6262/n1688 , \DP_OP_158_296_6262/n1670 ,
         \DP_OP_158_296_6262/n1663 , \DP_OP_158_296_6262/n1661 ,
         \DP_OP_158_296_6262/n1659 , \DP_OP_158_296_6262/n1656 ,
         \DP_OP_158_296_6262/n1647 , \DP_OP_158_296_6262/n1645 ,
         \DP_OP_158_296_6262/n1638 , \DP_OP_158_296_6262/n1627 ,
         \DP_OP_158_296_6262/n1625 , \DP_OP_158_296_6262/n1623 ,
         \DP_OP_158_296_6262/n1621 , \DP_OP_158_296_6262/n1618 ,
         \DP_OP_158_296_6262/n1607 , \DP_OP_158_296_6262/n1605 ,
         \DP_OP_158_296_6262/n1596 , \DP_OP_158_296_6262/n1583 ,
         \DP_OP_158_296_6262/n1581 , \DP_OP_158_296_6262/n1579 ,
         \DP_OP_158_296_6262/n1571 , \DP_OP_158_296_6262/n1558 ,
         \DP_OP_158_296_6262/n1556 , \DP_OP_158_296_6262/n1543 ,
         \DP_OP_158_296_6262/n1526 , \DP_OP_158_296_6262/n1524 ,
         \DP_OP_158_296_6262/n1522 , \DP_OP_158_296_6262/n1520 ,
         \DP_OP_158_296_6262/n1518 , \DP_OP_158_296_6262/n1515 ,
         \DP_OP_158_296_6262/n1502 , \DP_OP_158_296_6262/n1500 ,
         \DP_OP_158_296_6262/n1489 , \DP_OP_158_296_6262/n1474 ,
         \DP_OP_158_296_6262/n1472 , \DP_OP_158_296_6262/n1470 ,
         \DP_OP_158_296_6262/n1460 , \DP_OP_158_296_6262/n1445 ,
         \DP_OP_158_296_6262/n1443 , \DP_OP_158_296_6262/n1428 ,
         \DP_OP_158_296_6262/n1409 , \DP_OP_158_296_6262/n1407 ,
         \DP_OP_158_296_6262/n1405 , \DP_OP_158_296_6262/n1403 ,
         \DP_OP_158_296_6262/n1395 , \DP_OP_158_296_6262/n1380 ,
         \DP_OP_158_296_6262/n1378 , \DP_OP_158_296_6262/n1359 ,
         \DP_OP_158_296_6262/n1346 , \DP_OP_158_296_6262/n1344 ,
         \DP_OP_158_296_6262/n1342 , \DP_OP_158_296_6262/n1923 ,
         \DP_OP_158_296_6262/n1986 , \DP_OP_158_296_6262/n1933 ,
         \DP_OP_158_296_6262/n1932 , \DP_OP_158_296_6262/n1931 ,
         \DP_OP_158_296_6262/n1988 , \addr_calc/fft_write_calc/counter/N61 ,
         \DP_OP_158_296_6262/n822 , \DP_OP_158_296_6262/n820 ,
         \DP_OP_158_296_6262/n818 , \DP_OP_158_296_6262/n812 ,
         \DP_OP_158_296_6262/n796 , \DP_OP_158_296_6262/n794 ,
         \DP_OP_158_296_6262/n776 , \DP_OP_158_296_6262/n769 ,
         \DP_OP_158_296_6262/n767 , \DP_OP_158_296_6262/n765 ,
         \DP_OP_158_296_6262/n762 , \DP_OP_158_296_6262/n753 ,
         \DP_OP_158_296_6262/n751 , \DP_OP_158_296_6262/n744 ,
         \DP_OP_158_296_6262/n733 , \DP_OP_158_296_6262/n731 ,
         \DP_OP_158_296_6262/n729 , \DP_OP_158_296_6262/n727 ,
         \DP_OP_158_296_6262/n724 , \DP_OP_158_296_6262/n713 ,
         \DP_OP_158_296_6262/n711 , \DP_OP_158_296_6262/n702 ,
         \DP_OP_158_296_6262/n689 , \DP_OP_158_296_6262/n687 ,
         \DP_OP_158_296_6262/n685 , \DP_OP_158_296_6262/n677 ,
         \DP_OP_158_296_6262/n664 , \DP_OP_158_296_6262/n662 ,
         \DP_OP_158_296_6262/n649 , \DP_OP_158_296_6262/n632 ,
         \DP_OP_158_296_6262/n630 , \DP_OP_158_296_6262/n628 ,
         \DP_OP_158_296_6262/n626 , \DP_OP_158_296_6262/n621 ,
         \DP_OP_158_296_6262/n608 , \DP_OP_158_296_6262/n606 ,
         \DP_OP_158_296_6262/n595 , \DP_OP_158_296_6262/n580 ,
         \DP_OP_158_296_6262/n578 , \DP_OP_158_296_6262/n576 ,
         \DP_OP_158_296_6262/n566 , \DP_OP_158_296_6262/n549 ,
         \DP_OP_158_296_6262/n534 , \DP_OP_158_296_6262/n515 ,
         \DP_OP_158_296_6262/n513 , \DP_OP_158_296_6262/n511 ,
         \DP_OP_158_296_6262/n509 , \DP_OP_158_296_6262/n501 ,
         \DP_OP_158_296_6262/n486 , \DP_OP_158_296_6262/n484 ,
         \DP_OP_158_296_6262/n465 , \DP_OP_158_296_6262/n452 ,
         \DP_OP_158_296_6262/n450 , \DP_OP_158_296_6262/n1889 ,
         \DP_OP_158_296_6262/n1888 , \DP_OP_159_297_3515/n1014 ,
         \addr_calc/iir_read_calc/counter/N47 ,
         \addr_calc/iir_read_calc/counter/N49 ,
         \addr_calc/fir_write_calc/counter/N58 , \add_x_22_3/n65 ,
         \add_x_19_2/n50 , \add_x_19_2/n4 , \add_x_19_2/n195 , \add_x_19_2/n7 ,
         \add_x_19_2/n65 , \add_x_19_2/n198 , \add_x_19_2/n71 ,
         \add_x_19_2/n70 , \add_x_19_2/n119 , \add_x_19_2/n117 ,
         \add_x_19_2/n115 , \add_x_19_2/n114 , \add_x_19_2/n161 ,
         \add_x_19_2/n159 , \add_x_19_2/n158 ,
         \addr_calc/fir_read_calc/counter/N58 , \add_x_22_2/n65 ,
         \addr_calc/iir_write_calc/counter/N63 , \add_x_19_1/n99 ,
         \add_x_19_1/n204 , \add_x_19_1/n13 ,
         \addr_calc/fft_write_calc/counter/N69 , \add_x_19_1/n119 ,
         \add_x_19_1/n117 , \add_x_19_1/n115 , \add_x_19_1/n114 ,
         \add_x_19_1/n161 , \add_x_19_1/n159 , \add_x_19_1/n158 ,
         \add_x_19_1/n83 , \add_x_19_1/n157 , \add_x_19_1/n169 ,
         \add_x_19_1/n92 , \add_x_19_1/n113 , \add_x_19_1/n171 , n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2065, n2066, n2067, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813;

  NOR4XLTS U71 ( .A(n1785), .B(n1911), .C(\addr_calc/iir_read_calc/count[10] ), 
        .D(n2580), .Y(n816) );
  NOR4XLTS U197 ( .A(n1941), .B(\addr_calc/fft_write_calc/count[19] ), .C(
        n2020), .D(n1924), .Y(n846) );
  NOR4XLTS U274 ( .A(n2000), .B(n1877), .C(
        \addr_calc/fir_write_calc/count[10] ), .D(n1986), .Y(n867) );
  NOR4XLTS U288 ( .A(\addr_calc/fir_read_calc/count[16] ), .B(
        \addr_calc/fir_read_calc/count[15] ), .C(
        \addr_calc/fir_read_calc/count[14] ), .D(
        \addr_calc/fir_read_calc/count[13] ), .Y(n883) );
  NOR4XLTS U289 ( .A(n1994), .B(n1895), .C(\addr_calc/fir_read_calc/count[10] ), .D(n2007), .Y(n882) );
  NOR4XLTS U291 ( .A(\addr_calc/fir_read_calc/count[1] ), .B(
        \addr_calc/fir_read_calc/count[19] ), .C(n1988), .D(
        \addr_calc/fir_read_calc/count[17] ), .Y(n880) );
  NAND3X1TS U294 ( .A(n2055), .B(n2067), .C(n886), .Y(n885) );
  NAND3BX1TS U299 ( .AN(n884), .B(fir_write_done), .C(fir_read_done), .Y(n897)
         );
  OAI33XLTS U306 ( .A0(n891), .A1(n901), .A2(n1861), .B0(n899), .B1(n869), 
        .B2(iir_write_done), .Y(n1135) );
  NAND2X1TS U310 ( .A(n902), .B(n2311), .Y(n870) );
  NAND2X1TS U313 ( .A(n2336), .B(n872), .Y(n899) );
  NAND3X1TS U315 ( .A(n904), .B(n905), .C(n906), .Y(n903) );
  NAND3BX1TS U323 ( .AN(instruction[9]), .B(n2310), .C(
        \pla_top/instruction_valid ), .Y(n907) );
  NOR4XLTS U338 ( .A(n2044), .B(n1942), .C(n1940), .D(n2578), .Y(n921) );
  OA21XLTS U343 ( .A0(n796), .A1(n923), .B0(iir_get_req_reg), .Y(iir_get_req)
         );
  OA21XLTS U350 ( .A0(n798), .A1(n927), .B0(fir_get_req_reg), .Y(fir_get_req)
         );
  NOR4XLTS U365 ( .A(n2323), .B(n2327), .C(n933), .D(n932), .Y(
        \data_cntl/N256 ) );
  NOR4XLTS U371 ( .A(n2313), .B(n2315), .C(n937), .D(n1830), .Y(
        \data_cntl/N253 ) );
  NAND3X1TS U381 ( .A(n2815), .B(n2059), .C(n2586), .Y(n932) );
  TLATXLTS \data_cntl/fft_get_req_reg  ( .G(\data_cntl/N260 ), .D(
        \data_cntl/N261 ), .QN(n929) );
  TLATXLTS \data_cntl/fft_put_req_reg  ( .G(\data_cntl/N260 ), .D(
        \data_cntl/N259 ), .Q(fft_put_req_reg) );
  TLATXLTS \data_cntl/fir_put_req_reg  ( .G(\data_cntl/N263 ), .D(
        \data_cntl/N262 ), .Q(fir_put_req_reg) );
  TLATXLTS \data_cntl/iir_put_req_reg  ( .G(\data_cntl/N266 ), .D(
        \data_cntl/N265 ), .Q(iir_put_req_reg) );
  TLATXLTS \data_cntl/iir_get_req_reg  ( .G(\data_cntl/N266 ), .D(
        \data_cntl/N267 ), .Q(iir_get_req_reg) );
  TLATXLTS \data_cntl/fir_get_req_reg  ( .G(\data_cntl/N263 ), .D(
        \data_cntl/N264 ), .Q(fir_get_req_reg) );
  TLATXLTS \data_cntl/data_to_fft_reg  ( .G(\data_cntl/N250 ), .D(
        \data_cntl/N251 ), .Q(data_to_fft), .QN(\data_cntl/N63 ) );
  TLATXLTS \data_cntl/data_to_fir_reg  ( .G(\data_cntl/N255 ), .D(
        \data_cntl/N253 ), .Q(data_to_fir), .QN(\data_cntl/N99 ) );
  TLATXLTS \data_cntl/data_to_iir_reg  ( .G(\data_cntl/N258 ), .D(
        \data_cntl/N256 ), .Q(data_to_iir), .QN(\data_cntl/N191 ) );
  TLATXLTS \data_cntl/data_from_fft_reg  ( .G(\data_cntl/N250 ), .D(
        \data_cntl/N252 ), .Q(data_from_fft), .QN(\data_cntl/N9 ) );
  TLATXLTS \data_cntl/data_from_fir_reg  ( .G(\data_cntl/N255 ), .D(
        \data_cntl/N254 ), .Q(data_from_fir), .QN(\data_cntl/N95 ) );
  TLATXLTS \data_cntl/data_from_iir_reg  ( .G(\data_cntl/N258 ), .D(
        \data_cntl/N257 ), .Q(data_from_iir), .QN(\data_cntl/N159 ) );
  TLATXLTS \addr_calc/from_fir_go_reg  ( .G(\addr_calc/N220 ), .D(
        \data_cntl/N264 ), .Q(n2643), .QN(\addr_calc/N99 ) );
  TLATXLTS \addr_calc/to_fir_go_reg  ( .G(\addr_calc/N220 ), .D(
        \addr_calc/N219 ), .Q(n2644), .QN(\addr_calc/N95 ) );
  TLATXLTS \addr_calc/from_fft_go_reg  ( .G(\addr_calc/N216 ), .D(
        \data_cntl/N261 ), .Q(n2645), .QN(\addr_calc/N63 ) );
  TLATXLTS \addr_calc/to_fft_go_reg  ( .G(\addr_calc/N216 ), .D(
        \addr_calc/N217 ), .Q(n2646), .QN(\addr_calc/N9 ) );
  TLATXLTS \addr_calc/to_iir_go_reg  ( .G(\addr_calc/N224 ), .D(
        \addr_calc/N223 ), .Q(n2642), .QN(\addr_calc/N159 ) );
  TLATXLTS \addr_calc/from_iir_go_reg  ( .G(\addr_calc/N224 ), .D(
        \data_cntl/N267 ), .Q(n2641), .QN(\addr_calc/N191 ) );
  DFFQX1TS \pla_top/acc_done_reg  ( .D(n1134), .CK(clk), .Q(acc_done) );
  TBUFX2TS \data_cntl/fft_data_out_tri[31]  ( .A(n2360), .OE(n2690), .Y(
        fft_data_out[31]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[30]  ( .A(n2502), .OE(n2690), .Y(
        fft_data_out[30]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[29]  ( .A(n2518), .OE(n2690), .Y(
        fft_data_out[29]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[28]  ( .A(n2534), .OE(n2690), .Y(
        fft_data_out[28]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[27]  ( .A(n2356), .OE(n2691), .Y(
        fft_data_out[27]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[26]  ( .A(n2504), .OE(n2691), .Y(
        fft_data_out[26]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[25]  ( .A(n2520), .OE(n2691), .Y(
        fft_data_out[25]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[24]  ( .A(n2536), .OE(n2691), .Y(
        fft_data_out[24]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[23]  ( .A(n2352), .OE(n2692), .Y(
        fft_data_out[23]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[22]  ( .A(n2506), .OE(n2692), .Y(
        fft_data_out[22]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[21]  ( .A(n2522), .OE(n2692), .Y(
        fft_data_out[21]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[20]  ( .A(n2538), .OE(n2692), .Y(
        fft_data_out[20]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[19]  ( .A(n2348), .OE(n2693), .Y(
        fft_data_out[19]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[18]  ( .A(n2508), .OE(n2693), .Y(
        fft_data_out[18]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[17]  ( .A(n2524), .OE(n2693), .Y(
        fft_data_out[17]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[16]  ( .A(n2540), .OE(n2693), .Y(
        fft_data_out[16]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[15]  ( .A(n2346), .OE(n2694), .Y(
        fft_data_out[15]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[14]  ( .A(n2510), .OE(n2694), .Y(
        fft_data_out[14]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[13]  ( .A(n2526), .OE(n2694), .Y(
        fft_data_out[13]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[12]  ( .A(n2542), .OE(n2694), .Y(
        fft_data_out[12]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[11]  ( .A(n2350), .OE(n2695), .Y(
        fft_data_out[11]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[10]  ( .A(n2512), .OE(n2695), .Y(
        fft_data_out[10]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[9]  ( .A(n2528), .OE(n2695), .Y(
        fft_data_out[9]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[8]  ( .A(n2544), .OE(n2695), .Y(
        fft_data_out[8]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[7]  ( .A(n2354), .OE(n2696), .Y(
        fft_data_out[7]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[6]  ( .A(n2514), .OE(n2696), .Y(
        fft_data_out[6]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[5]  ( .A(n2530), .OE(n2696), .Y(
        fft_data_out[5]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[4]  ( .A(n2546), .OE(n2696), .Y(
        fft_data_out[4]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[3]  ( .A(n2358), .OE(n2697), .Y(
        fft_data_out[3]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[2]  ( .A(n2516), .OE(n2697), .Y(
        fft_data_out[2]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[1]  ( .A(n2532), .OE(n2697), .Y(
        fft_data_out[1]) );
  TBUFX2TS \data_cntl/fft_data_out_tri[0]  ( .A(n2548), .OE(n2697), .Y(
        fft_data_out[0]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[31]  ( .A(n2360), .OE(n2708), .Y(
        fir_data_out[31]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[30]  ( .A(n2502), .OE(n2708), .Y(
        fir_data_out[30]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[29]  ( .A(n2518), .OE(n2708), .Y(
        fir_data_out[29]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[28]  ( .A(n2534), .OE(n2708), .Y(
        fir_data_out[28]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[27]  ( .A(n2356), .OE(n2709), .Y(
        fir_data_out[27]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[26]  ( .A(n2504), .OE(n2709), .Y(
        fir_data_out[26]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[25]  ( .A(n2520), .OE(n2709), .Y(
        fir_data_out[25]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[24]  ( .A(n2536), .OE(n2709), .Y(
        fir_data_out[24]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[23]  ( .A(n2352), .OE(n2710), .Y(
        fir_data_out[23]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[22]  ( .A(n2506), .OE(n2710), .Y(
        fir_data_out[22]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[21]  ( .A(n2522), .OE(n2710), .Y(
        fir_data_out[21]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[20]  ( .A(n2538), .OE(n2710), .Y(
        fir_data_out[20]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[19]  ( .A(n2348), .OE(n2711), .Y(
        fir_data_out[19]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[18]  ( .A(n2508), .OE(n2711), .Y(
        fir_data_out[18]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[17]  ( .A(n2524), .OE(n2711), .Y(
        fir_data_out[17]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[16]  ( .A(n2540), .OE(n2711), .Y(
        fir_data_out[16]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[15]  ( .A(n2346), .OE(n2712), .Y(
        fir_data_out[15]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[14]  ( .A(n2510), .OE(n2712), .Y(
        fir_data_out[14]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[13]  ( .A(n2526), .OE(n2712), .Y(
        fir_data_out[13]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[12]  ( .A(n2542), .OE(n2712), .Y(
        fir_data_out[12]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[11]  ( .A(n2350), .OE(n2713), .Y(
        fir_data_out[11]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[10]  ( .A(n2512), .OE(n2713), .Y(
        fir_data_out[10]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[9]  ( .A(n2528), .OE(n2713), .Y(
        fir_data_out[9]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[8]  ( .A(n2544), .OE(n2713), .Y(
        fir_data_out[8]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[7]  ( .A(n2354), .OE(n2714), .Y(
        fir_data_out[7]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[6]  ( .A(n2514), .OE(n2714), .Y(
        fir_data_out[6]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[5]  ( .A(n2530), .OE(n2714), .Y(
        fir_data_out[5]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[4]  ( .A(n2546), .OE(n2714), .Y(
        fir_data_out[4]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[3]  ( .A(n2358), .OE(n2715), .Y(
        fir_data_out[3]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[2]  ( .A(n2516), .OE(n2715), .Y(
        fir_data_out[2]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[1]  ( .A(n2532), .OE(n2715), .Y(
        fir_data_out[1]) );
  TBUFX2TS \data_cntl/fir_data_out_tri[0]  ( .A(n2548), .OE(n2715), .Y(
        fir_data_out[0]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[31]  ( .A(n2360), .OE(n2726), .Y(
        iir_data_out[31]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[30]  ( .A(n2502), .OE(n2726), .Y(
        iir_data_out[30]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[29]  ( .A(n2518), .OE(n2726), .Y(
        iir_data_out[29]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[28]  ( .A(n2534), .OE(n2726), .Y(
        iir_data_out[28]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[27]  ( .A(n2356), .OE(n2727), .Y(
        iir_data_out[27]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[26]  ( .A(n2504), .OE(n2727), .Y(
        iir_data_out[26]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[25]  ( .A(n2520), .OE(n2727), .Y(
        iir_data_out[25]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[24]  ( .A(n2536), .OE(n2727), .Y(
        iir_data_out[24]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[23]  ( .A(n2352), .OE(n2728), .Y(
        iir_data_out[23]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[22]  ( .A(n2506), .OE(n2728), .Y(
        iir_data_out[22]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[21]  ( .A(n2522), .OE(n2728), .Y(
        iir_data_out[21]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[20]  ( .A(n2538), .OE(n2728), .Y(
        iir_data_out[20]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[19]  ( .A(n2348), .OE(n2729), .Y(
        iir_data_out[19]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[18]  ( .A(n2508), .OE(n2729), .Y(
        iir_data_out[18]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[17]  ( .A(n2524), .OE(n2729), .Y(
        iir_data_out[17]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[16]  ( .A(n2540), .OE(n2729), .Y(
        iir_data_out[16]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[15]  ( .A(n2346), .OE(n2730), .Y(
        iir_data_out[15]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[14]  ( .A(n2510), .OE(n2730), .Y(
        iir_data_out[14]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[13]  ( .A(n2526), .OE(n2730), .Y(
        iir_data_out[13]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[12]  ( .A(n2542), .OE(n2730), .Y(
        iir_data_out[12]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[11]  ( .A(n2350), .OE(n2731), .Y(
        iir_data_out[11]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[10]  ( .A(n2512), .OE(n2731), .Y(
        iir_data_out[10]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[9]  ( .A(n2528), .OE(n2731), .Y(
        iir_data_out[9]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[8]  ( .A(n2544), .OE(n2731), .Y(
        iir_data_out[8]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[7]  ( .A(n2354), .OE(n2732), .Y(
        iir_data_out[7]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[6]  ( .A(n2514), .OE(n2732), .Y(
        iir_data_out[6]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[5]  ( .A(n2530), .OE(n2732), .Y(
        iir_data_out[5]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[4]  ( .A(n2546), .OE(n2732), .Y(
        iir_data_out[4]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[3]  ( .A(n2358), .OE(n2733), .Y(
        iir_data_out[3]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[2]  ( .A(n2516), .OE(n2733), .Y(
        iir_data_out[2]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[1]  ( .A(n2532), .OE(n2733), .Y(
        iir_data_out[1]) );
  TBUFX2TS \data_cntl/iir_data_out_tri[0]  ( .A(n2548), .OE(n2733), .Y(
        iir_data_out[0]) );
  TBUFX2TS \data_cntl/data_bus_tri[31]  ( .A(n2308), .OE(n2681), .Y(
        data_bus[31]) );
  TBUFX2TS \data_cntl/data_bus_tri[30]  ( .A(n2304), .OE(n2681), .Y(
        data_bus[30]) );
  TBUFX2TS \data_cntl/data_bus_tri[29]  ( .A(n2300), .OE(n2681), .Y(
        data_bus[29]) );
  TBUFX2TS \data_cntl/data_bus_tri[28]  ( .A(n2296), .OE(n2681), .Y(
        data_bus[28]) );
  TBUFX2TS \data_cntl/data_bus_tri[27]  ( .A(n2292), .OE(n2682), .Y(
        data_bus[27]) );
  TBUFX2TS \data_cntl/data_bus_tri[26]  ( .A(n2288), .OE(n2682), .Y(
        data_bus[26]) );
  TBUFX2TS \data_cntl/data_bus_tri[25]  ( .A(n2284), .OE(n2682), .Y(
        data_bus[25]) );
  TBUFX2TS \data_cntl/data_bus_tri[24]  ( .A(n2280), .OE(n2682), .Y(
        data_bus[24]) );
  TBUFX2TS \data_cntl/data_bus_tri[23]  ( .A(n2276), .OE(n2683), .Y(
        data_bus[23]) );
  TBUFX2TS \data_cntl/data_bus_tri[22]  ( .A(n2272), .OE(n2683), .Y(
        data_bus[22]) );
  TBUFX2TS \data_cntl/data_bus_tri[21]  ( .A(n2268), .OE(n2683), .Y(
        data_bus[21]) );
  TBUFX2TS \data_cntl/data_bus_tri[20]  ( .A(n2264), .OE(n2683), .Y(
        data_bus[20]) );
  TBUFX2TS \data_cntl/data_bus_tri[19]  ( .A(n2260), .OE(n2684), .Y(
        data_bus[19]) );
  TBUFX2TS \data_cntl/data_bus_tri[18]  ( .A(n2256), .OE(n2684), .Y(
        data_bus[18]) );
  TBUFX2TS \data_cntl/data_bus_tri[17]  ( .A(n2252), .OE(n2684), .Y(
        data_bus[17]) );
  TBUFX2TS \data_cntl/data_bus_tri[16]  ( .A(n2248), .OE(n2684), .Y(
        data_bus[16]) );
  TBUFX2TS \data_cntl/data_bus_tri[15]  ( .A(n2244), .OE(n2685), .Y(
        data_bus[15]) );
  TBUFX2TS \data_cntl/data_bus_tri[14]  ( .A(n2240), .OE(n2685), .Y(
        data_bus[14]) );
  TBUFX2TS \data_cntl/data_bus_tri[13]  ( .A(n2236), .OE(n2685), .Y(
        data_bus[13]) );
  TBUFX2TS \data_cntl/data_bus_tri[12]  ( .A(n2232), .OE(n2685), .Y(
        data_bus[12]) );
  TBUFX2TS \data_cntl/data_bus_tri[11]  ( .A(n2228), .OE(n2686), .Y(
        data_bus[11]) );
  TBUFX2TS \data_cntl/data_bus_tri[10]  ( .A(n2224), .OE(n2686), .Y(
        data_bus[10]) );
  TBUFX2TS \data_cntl/data_bus_tri[9]  ( .A(n2220), .OE(n2686), .Y(data_bus[9]) );
  TBUFX2TS \data_cntl/data_bus_tri[8]  ( .A(n2216), .OE(n2686), .Y(data_bus[8]) );
  TBUFX2TS \data_cntl/data_bus_tri[7]  ( .A(n2212), .OE(n2687), .Y(data_bus[7]) );
  TBUFX2TS \data_cntl/data_bus_tri[6]  ( .A(n2208), .OE(n2687), .Y(data_bus[6]) );
  TBUFX2TS \data_cntl/data_bus_tri[5]  ( .A(n2204), .OE(n2687), .Y(data_bus[5]) );
  TBUFX2TS \data_cntl/data_bus_tri[4]  ( .A(n2200), .OE(n2687), .Y(data_bus[4]) );
  TBUFX2TS \data_cntl/data_bus_tri[3]  ( .A(n2196), .OE(n2688), .Y(data_bus[3]) );
  TBUFX2TS \data_cntl/data_bus_tri[2]  ( .A(n2192), .OE(n2688), .Y(data_bus[2]) );
  TBUFX2TS \data_cntl/data_bus_tri[1]  ( .A(n2188), .OE(n2688), .Y(data_bus[1]) );
  TBUFX2TS \data_cntl/data_bus_tri[0]  ( .A(n2184), .OE(n2688), .Y(data_bus[0]) );
  TBUFX2TS \data_cntl/data_bus_tri2[31]  ( .A(n2180), .OE(n2699), .Y(
        data_bus[31]) );
  TBUFX2TS \data_cntl/data_bus_tri2[30]  ( .A(n2176), .OE(n2699), .Y(
        data_bus[30]) );
  TBUFX2TS \data_cntl/data_bus_tri2[29]  ( .A(n2172), .OE(n2699), .Y(
        data_bus[29]) );
  TBUFX2TS \data_cntl/data_bus_tri2[28]  ( .A(n2168), .OE(n2699), .Y(
        data_bus[28]) );
  TBUFX2TS \data_cntl/data_bus_tri2[27]  ( .A(n2164), .OE(n2700), .Y(
        data_bus[27]) );
  TBUFX2TS \data_cntl/data_bus_tri2[26]  ( .A(n2160), .OE(n2700), .Y(
        data_bus[26]) );
  TBUFX2TS \data_cntl/data_bus_tri2[25]  ( .A(n2156), .OE(n2700), .Y(
        data_bus[25]) );
  TBUFX2TS \data_cntl/data_bus_tri2[24]  ( .A(n2152), .OE(n2700), .Y(
        data_bus[24]) );
  TBUFX2TS \data_cntl/data_bus_tri2[23]  ( .A(n2148), .OE(n2701), .Y(
        data_bus[23]) );
  TBUFX2TS \data_cntl/data_bus_tri2[22]  ( .A(n2144), .OE(n2701), .Y(
        data_bus[22]) );
  TBUFX2TS \data_cntl/data_bus_tri2[21]  ( .A(n2140), .OE(n2701), .Y(
        data_bus[21]) );
  TBUFX2TS \data_cntl/data_bus_tri2[20]  ( .A(n2136), .OE(n2701), .Y(
        data_bus[20]) );
  TBUFX2TS \data_cntl/data_bus_tri2[19]  ( .A(n2132), .OE(n2702), .Y(
        data_bus[19]) );
  TBUFX2TS \data_cntl/data_bus_tri2[18]  ( .A(n2128), .OE(n2702), .Y(
        data_bus[18]) );
  TBUFX2TS \data_cntl/data_bus_tri2[17]  ( .A(n2124), .OE(n2702), .Y(
        data_bus[17]) );
  TBUFX2TS \data_cntl/data_bus_tri2[16]  ( .A(n2120), .OE(n2702), .Y(
        data_bus[16]) );
  TBUFX2TS \data_cntl/data_bus_tri2[15]  ( .A(n2118), .OE(n2703), .Y(
        data_bus[15]) );
  TBUFX2TS \data_cntl/data_bus_tri2[14]  ( .A(n2122), .OE(n2703), .Y(
        data_bus[14]) );
  TBUFX2TS \data_cntl/data_bus_tri2[13]  ( .A(n2126), .OE(n2703), .Y(
        data_bus[13]) );
  TBUFX2TS \data_cntl/data_bus_tri2[12]  ( .A(n2130), .OE(n2703), .Y(
        data_bus[12]) );
  TBUFX2TS \data_cntl/data_bus_tri2[11]  ( .A(n2134), .OE(n2704), .Y(
        data_bus[11]) );
  TBUFX2TS \data_cntl/data_bus_tri2[10]  ( .A(n2138), .OE(n2704), .Y(
        data_bus[10]) );
  TBUFX2TS \data_cntl/data_bus_tri2[9]  ( .A(n2142), .OE(n2704), .Y(
        data_bus[9]) );
  TBUFX2TS \data_cntl/data_bus_tri2[8]  ( .A(n2146), .OE(n2704), .Y(
        data_bus[8]) );
  TBUFX2TS \data_cntl/data_bus_tri2[7]  ( .A(n2150), .OE(n2705), .Y(
        data_bus[7]) );
  TBUFX2TS \data_cntl/data_bus_tri2[6]  ( .A(n2154), .OE(n2705), .Y(
        data_bus[6]) );
  TBUFX2TS \data_cntl/data_bus_tri2[5]  ( .A(n2158), .OE(n2705), .Y(
        data_bus[5]) );
  TBUFX2TS \data_cntl/data_bus_tri2[4]  ( .A(n2162), .OE(n2705), .Y(
        data_bus[4]) );
  TBUFX2TS \data_cntl/data_bus_tri2[3]  ( .A(n2166), .OE(n2706), .Y(
        data_bus[3]) );
  TBUFX2TS \data_cntl/data_bus_tri2[2]  ( .A(n2170), .OE(n2706), .Y(
        data_bus[2]) );
  TBUFX2TS \data_cntl/data_bus_tri2[1]  ( .A(n2174), .OE(n2706), .Y(
        data_bus[1]) );
  TBUFX2TS \data_cntl/data_bus_tri2[0]  ( .A(n2178), .OE(n2706), .Y(
        data_bus[0]) );
  TBUFX2TS \data_cntl/data_bus_tri3[31]  ( .A(n2182), .OE(n2717), .Y(
        data_bus[31]) );
  TBUFX2TS \data_cntl/data_bus_tri3[30]  ( .A(n2186), .OE(n2717), .Y(
        data_bus[30]) );
  TBUFX2TS \data_cntl/data_bus_tri3[29]  ( .A(n2190), .OE(n2717), .Y(
        data_bus[29]) );
  TBUFX2TS \data_cntl/data_bus_tri3[28]  ( .A(n2194), .OE(n2717), .Y(
        data_bus[28]) );
  TBUFX2TS \data_cntl/data_bus_tri3[27]  ( .A(n2198), .OE(n2718), .Y(
        data_bus[27]) );
  TBUFX2TS \data_cntl/data_bus_tri3[26]  ( .A(n2202), .OE(n2718), .Y(
        data_bus[26]) );
  TBUFX2TS \data_cntl/data_bus_tri3[25]  ( .A(n2206), .OE(n2718), .Y(
        data_bus[25]) );
  TBUFX2TS \data_cntl/data_bus_tri3[24]  ( .A(n2210), .OE(n2718), .Y(
        data_bus[24]) );
  TBUFX2TS \data_cntl/data_bus_tri3[23]  ( .A(n2214), .OE(n2719), .Y(
        data_bus[23]) );
  TBUFX2TS \data_cntl/data_bus_tri3[22]  ( .A(n2218), .OE(n2719), .Y(
        data_bus[22]) );
  TBUFX2TS \data_cntl/data_bus_tri3[21]  ( .A(n2222), .OE(n2719), .Y(
        data_bus[21]) );
  TBUFX2TS \data_cntl/data_bus_tri3[20]  ( .A(n2226), .OE(n2719), .Y(
        data_bus[20]) );
  TBUFX2TS \data_cntl/data_bus_tri3[19]  ( .A(n2230), .OE(n2720), .Y(
        data_bus[19]) );
  TBUFX2TS \data_cntl/data_bus_tri3[18]  ( .A(n2234), .OE(n2720), .Y(
        data_bus[18]) );
  TBUFX2TS \data_cntl/data_bus_tri3[17]  ( .A(n2238), .OE(n2720), .Y(
        data_bus[17]) );
  TBUFX2TS \data_cntl/data_bus_tri3[16]  ( .A(n2242), .OE(n2720), .Y(
        data_bus[16]) );
  TBUFX2TS \data_cntl/data_bus_tri3[15]  ( .A(n2246), .OE(n2721), .Y(
        data_bus[15]) );
  TBUFX2TS \data_cntl/data_bus_tri3[14]  ( .A(n2250), .OE(n2721), .Y(
        data_bus[14]) );
  TBUFX2TS \data_cntl/data_bus_tri3[13]  ( .A(n2254), .OE(n2721), .Y(
        data_bus[13]) );
  TBUFX2TS \data_cntl/data_bus_tri3[12]  ( .A(n2258), .OE(n2721), .Y(
        data_bus[12]) );
  TBUFX2TS \data_cntl/data_bus_tri3[11]  ( .A(n2262), .OE(n2722), .Y(
        data_bus[11]) );
  TBUFX2TS \data_cntl/data_bus_tri3[10]  ( .A(n2266), .OE(n2722), .Y(
        data_bus[10]) );
  TBUFX2TS \data_cntl/data_bus_tri3[9]  ( .A(n2270), .OE(n2722), .Y(
        data_bus[9]) );
  TBUFX2TS \data_cntl/data_bus_tri3[8]  ( .A(n2274), .OE(n2722), .Y(
        data_bus[8]) );
  TBUFX2TS \data_cntl/data_bus_tri3[7]  ( .A(n2278), .OE(n2723), .Y(
        data_bus[7]) );
  TBUFX2TS \data_cntl/data_bus_tri3[6]  ( .A(n2282), .OE(n2723), .Y(
        data_bus[6]) );
  TBUFX2TS \data_cntl/data_bus_tri3[5]  ( .A(n2286), .OE(n2723), .Y(
        data_bus[5]) );
  TBUFX2TS \data_cntl/data_bus_tri3[4]  ( .A(n2290), .OE(n2723), .Y(
        data_bus[4]) );
  TBUFX2TS \data_cntl/data_bus_tri3[3]  ( .A(n2294), .OE(n2724), .Y(
        data_bus[3]) );
  TBUFX2TS \data_cntl/data_bus_tri3[2]  ( .A(n2298), .OE(n2724), .Y(
        data_bus[2]) );
  TBUFX2TS \data_cntl/data_bus_tri3[1]  ( .A(n2302), .OE(n2724), .Y(
        data_bus[1]) );
  TBUFX2TS \data_cntl/data_bus_tri3[0]  ( .A(n2306), .OE(n2724), .Y(
        data_bus[0]) );
  TBUFX2TS \addr_calc/addr_tri[0]  ( .A(\addr_calc/fft_read_addr[0] ), .OE(
        n2742), .Y(addr[0]) );
  TBUFX2TS \addr_calc/addr_tri2[0]  ( .A(\addr_calc/fft_write_addr[0] ), .OE(
        n2750), .Y(addr[0]) );
  TBUFX2TS \addr_calc/addr_tri3[0]  ( .A(\addr_calc/fir_read_addr[0] ), .OE(
        n2758), .Y(addr[0]) );
  TBUFX2TS \addr_calc/addr_tri4[0]  ( .A(\addr_calc/fir_write_addr[0] ), .OE(
        n2766), .Y(addr[0]) );
  TBUFX2TS \addr_calc/addr_tri5[0]  ( .A(\addr_calc/iir_read_addr[0] ), .OE(
        n2774), .Y(addr[0]) );
  TBUFX2TS \addr_calc/addr_tri6[0]  ( .A(\addr_calc/iir_write_addr[0] ), .OE(
        n2782), .Y(addr[0]) );
  TBUFX2TS \addr_calc/addr_tri[3]  ( .A(\addr_calc/fft_read_addr[3] ), .OE(
        n2742), .Y(addr[3]) );
  TBUFX2TS \addr_calc/addr_tri2[4]  ( .A(\addr_calc/fft_write_addr[4] ), .OE(
        n2749), .Y(addr[4]) );
  TBUFX2TS \addr_calc/addr_tri2[3]  ( .A(\addr_calc/fft_write_addr[3] ), .OE(
        n2750), .Y(addr[3]) );
  TBUFX2TS \addr_calc/addr_tri3[4]  ( .A(\addr_calc/fir_read_addr[4] ), .OE(
        n2757), .Y(addr[4]) );
  TBUFX2TS \addr_calc/addr_tri3[3]  ( .A(\addr_calc/fir_read_addr[3] ), .OE(
        n2758), .Y(addr[3]) );
  TBUFX2TS \addr_calc/addr_tri4[4]  ( .A(\addr_calc/fir_write_addr[4] ), .OE(
        n2765), .Y(addr[4]) );
  TBUFX2TS \addr_calc/addr_tri4[3]  ( .A(\addr_calc/fir_write_addr[3] ), .OE(
        n2766), .Y(addr[3]) );
  TBUFX2TS \addr_calc/addr_tri5[3]  ( .A(\addr_calc/iir_read_addr[3] ), .OE(
        n2774), .Y(addr[3]) );
  TBUFX2TS \addr_calc/addr_tri6[4]  ( .A(\addr_calc/iir_write_addr[4] ), .OE(
        n2781), .Y(addr[4]) );
  TBUFX2TS \addr_calc/addr_tri6[3]  ( .A(\addr_calc/iir_write_addr[3] ), .OE(
        n2782), .Y(addr[3]) );
  TBUFX2TS \addr_calc/addr_tri[1]  ( .A(\addr_calc/fft_read_addr[1] ), .OE(
        n2742), .Y(addr[1]) );
  TBUFX2TS \addr_calc/addr_tri2[2]  ( .A(\addr_calc/fft_write_addr[2] ), .OE(
        n2750), .Y(addr[2]) );
  TBUFX2TS \addr_calc/addr_tri2[1]  ( .A(\addr_calc/fft_write_addr[1] ), .OE(
        n2750), .Y(addr[1]) );
  TBUFX2TS \addr_calc/addr_tri3[2]  ( .A(\addr_calc/fir_read_addr[2] ), .OE(
        n2758), .Y(addr[2]) );
  TBUFX2TS \addr_calc/addr_tri3[1]  ( .A(\addr_calc/fir_read_addr[1] ), .OE(
        n2758), .Y(addr[1]) );
  TBUFX2TS \addr_calc/addr_tri4[2]  ( .A(\addr_calc/fir_write_addr[2] ), .OE(
        n2766), .Y(addr[2]) );
  TBUFX2TS \addr_calc/addr_tri4[1]  ( .A(\addr_calc/fir_write_addr[1] ), .OE(
        n2766), .Y(addr[1]) );
  TBUFX2TS \addr_calc/addr_tri5[1]  ( .A(\addr_calc/iir_read_addr[1] ), .OE(
        n2774), .Y(addr[1]) );
  TBUFX2TS \addr_calc/addr_tri6[2]  ( .A(\addr_calc/iir_write_addr[2] ), .OE(
        n2782), .Y(addr[2]) );
  TBUFX2TS \addr_calc/addr_tri6[1]  ( .A(\addr_calc/iir_write_addr[1] ), .OE(
        n2782), .Y(addr[1]) );
  DFFQX1TS \pla_top/instruction_valid_reg  ( .D(\pla_top/N59 ), .CK(clk), .Q(
        \pla_top/instruction_valid ) );
  DFFQX1TS \pla_top/iir_enable_reg  ( .D(n1135), .CK(clk), .Q(n2815) );
  TBUFX2TS \addr_calc/addr_tri[29]  ( .A(\addr_calc/fft_read_addr[29] ), .OE(
        n2735), .Y(addr[29]) );
  TBUFX2TS \addr_calc/addr_tri[16]  ( .A(\addr_calc/fft_read_addr[16] ), .OE(
        n2738), .Y(addr[16]) );
  TBUFX4TS \addr_calc/addr_tri[13]  ( .A(\addr_calc/fft_read_addr[13] ), .OE(
        n2739), .Y(addr[13]) );
  TBUFX2TS \addr_calc/addr_tri[10]  ( .A(\addr_calc/fft_read_addr[10] ), .OE(
        n2740), .Y(addr[10]) );
  TBUFX2TS \addr_calc/addr_tri[9]  ( .A(\addr_calc/fft_read_addr[9] ), .OE(
        n2740), .Y(addr[9]) );
  TBUFX2TS \addr_calc/addr_tri[7]  ( .A(\addr_calc/fft_read_addr[7] ), .OE(
        n2741), .Y(addr[7]) );
  TBUFX2TS \addr_calc/addr_tri[4]  ( .A(\addr_calc/fft_read_addr[4] ), .OE(
        n2741), .Y(addr[4]) );
  TBUFX2TS \addr_calc/addr_tri2[29]  ( .A(\addr_calc/fft_write_addr[29] ), 
        .OE(n2743), .Y(addr[29]) );
  TBUFX2TS \addr_calc/addr_tri2[16]  ( .A(\addr_calc/fft_write_addr[16] ), 
        .OE(n2746), .Y(addr[16]) );
  TBUFX2TS \addr_calc/addr_tri2[10]  ( .A(\addr_calc/fft_write_addr[10] ), 
        .OE(n2748), .Y(addr[10]) );
  TBUFX2TS \addr_calc/addr_tri2[9]  ( .A(\addr_calc/fft_write_addr[9] ), .OE(
        n2748), .Y(addr[9]) );
  TBUFX2TS \addr_calc/addr_tri2[7]  ( .A(\addr_calc/fft_write_addr[7] ), .OE(
        n2749), .Y(addr[7]) );
  TBUFX2TS \addr_calc/addr_tri3[29]  ( .A(\addr_calc/fir_read_addr[29] ), .OE(
        n2751), .Y(addr[29]) );
  TBUFX2TS \addr_calc/addr_tri3[16]  ( .A(\addr_calc/fir_read_addr[16] ), .OE(
        n2754), .Y(addr[16]) );
  TBUFX2TS \addr_calc/addr_tri3[10]  ( .A(\addr_calc/fir_read_addr[10] ), .OE(
        n2756), .Y(addr[10]) );
  TBUFX2TS \addr_calc/addr_tri3[9]  ( .A(\addr_calc/fir_read_addr[9] ), .OE(
        n2756), .Y(addr[9]) );
  TBUFX2TS \addr_calc/addr_tri3[7]  ( .A(\addr_calc/fir_read_addr[7] ), .OE(
        n2757), .Y(addr[7]) );
  TBUFX2TS \addr_calc/addr_tri4[29]  ( .A(\addr_calc/fir_write_addr[29] ), 
        .OE(n2759), .Y(addr[29]) );
  TBUFX2TS \addr_calc/addr_tri4[16]  ( .A(\addr_calc/fir_write_addr[16] ), 
        .OE(n2762), .Y(addr[16]) );
  TBUFX2TS \addr_calc/addr_tri4[10]  ( .A(\addr_calc/fir_write_addr[10] ), 
        .OE(n2764), .Y(addr[10]) );
  TBUFX2TS \addr_calc/addr_tri4[9]  ( .A(\addr_calc/fir_write_addr[9] ), .OE(
        n2764), .Y(addr[9]) );
  TBUFX2TS \addr_calc/addr_tri4[7]  ( .A(\addr_calc/fir_write_addr[7] ), .OE(
        n2765), .Y(addr[7]) );
  TBUFX2TS \addr_calc/addr_tri5[16]  ( .A(\addr_calc/iir_read_addr[16] ), .OE(
        n2770), .Y(addr[16]) );
  TBUFX2TS \addr_calc/addr_tri5[10]  ( .A(\addr_calc/iir_read_addr[10] ), .OE(
        n2772), .Y(addr[10]) );
  TBUFX2TS \addr_calc/addr_tri5[9]  ( .A(\addr_calc/iir_read_addr[9] ), .OE(
        n2772), .Y(addr[9]) );
  TBUFX2TS \addr_calc/addr_tri5[7]  ( .A(\addr_calc/iir_read_addr[7] ), .OE(
        n2773), .Y(addr[7]) );
  TBUFX2TS \addr_calc/addr_tri5[4]  ( .A(\addr_calc/iir_read_addr[4] ), .OE(
        n2773), .Y(addr[4]) );
  TBUFX2TS \addr_calc/addr_tri6[29]  ( .A(\addr_calc/iir_write_addr[29] ), 
        .OE(n2775), .Y(addr[29]) );
  TBUFX2TS \addr_calc/addr_tri6[16]  ( .A(\addr_calc/iir_write_addr[16] ), 
        .OE(n2778), .Y(addr[16]) );
  TBUFX2TS \addr_calc/addr_tri6[10]  ( .A(\addr_calc/iir_write_addr[10] ), 
        .OE(n2780), .Y(addr[10]) );
  TBUFX2TS \addr_calc/addr_tri6[9]  ( .A(\addr_calc/iir_write_addr[9] ), .OE(
        n2780), .Y(addr[9]) );
  TBUFX2TS \addr_calc/addr_tri6[7]  ( .A(\addr_calc/iir_write_addr[7] ), .OE(
        n2781), .Y(addr[7]) );
  TBUFX2TS \addr_calc/addr_tri[12]  ( .A(\addr_calc/fft_read_addr[12] ), .OE(
        n2739), .Y(addr[12]) );
  TBUFX2TS \addr_calc/addr_tri[11]  ( .A(\addr_calc/fft_read_addr[11] ), .OE(
        n2740), .Y(addr[11]) );
  TBUFX2TS \addr_calc/addr_tri[8]  ( .A(\addr_calc/fft_read_addr[8] ), .OE(
        n2740), .Y(addr[8]) );
  TBUFX2TS \addr_calc/addr_tri[6]  ( .A(\addr_calc/fft_read_addr[6] ), .OE(
        n2741), .Y(addr[6]) );
  TBUFX2TS \addr_calc/addr_tri[5]  ( .A(\addr_calc/fft_read_addr[5] ), .OE(
        n2741), .Y(addr[5]) );
  TBUFX2TS \addr_calc/addr_tri[2]  ( .A(\addr_calc/fft_read_addr[2] ), .OE(
        n2742), .Y(addr[2]) );
  TBUFX2TS \addr_calc/addr_tri2[24]  ( .A(\addr_calc/fft_write_addr[24] ), 
        .OE(n2744), .Y(addr[24]) );
  TBUFX2TS \addr_calc/addr_tri2[20]  ( .A(\addr_calc/fft_write_addr[20] ), 
        .OE(n2745), .Y(addr[20]) );
  TBUFX2TS \addr_calc/addr_tri2[12]  ( .A(\addr_calc/fft_write_addr[12] ), 
        .OE(n2747), .Y(addr[12]) );
  TBUFX2TS \addr_calc/addr_tri2[11]  ( .A(\addr_calc/fft_write_addr[11] ), 
        .OE(n2748), .Y(addr[11]) );
  TBUFX2TS \addr_calc/addr_tri2[8]  ( .A(\addr_calc/fft_write_addr[8] ), .OE(
        n2748), .Y(addr[8]) );
  TBUFX2TS \addr_calc/addr_tri2[6]  ( .A(\addr_calc/fft_write_addr[6] ), .OE(
        n2749), .Y(addr[6]) );
  TBUFX2TS \addr_calc/addr_tri2[5]  ( .A(\addr_calc/fft_write_addr[5] ), .OE(
        n2749), .Y(addr[5]) );
  TBUFX2TS \addr_calc/addr_tri3[24]  ( .A(\addr_calc/fir_read_addr[24] ), .OE(
        n2752), .Y(addr[24]) );
  TBUFX2TS \addr_calc/addr_tri3[14]  ( .A(\addr_calc/fir_read_addr[14] ), .OE(
        n2755), .Y(addr[14]) );
  TBUFX2TS \addr_calc/addr_tri3[12]  ( .A(\addr_calc/fir_read_addr[12] ), .OE(
        n2755), .Y(addr[12]) );
  TBUFX2TS \addr_calc/addr_tri3[11]  ( .A(\addr_calc/fir_read_addr[11] ), .OE(
        n2756), .Y(addr[11]) );
  TBUFX2TS \addr_calc/addr_tri3[8]  ( .A(\addr_calc/fir_read_addr[8] ), .OE(
        n2756), .Y(addr[8]) );
  TBUFX2TS \addr_calc/addr_tri3[6]  ( .A(\addr_calc/fir_read_addr[6] ), .OE(
        n2757), .Y(addr[6]) );
  TBUFX2TS \addr_calc/addr_tri3[5]  ( .A(\addr_calc/fir_read_addr[5] ), .OE(
        n2757), .Y(addr[5]) );
  TBUFX2TS \addr_calc/addr_tri4[24]  ( .A(\addr_calc/fir_write_addr[24] ), 
        .OE(n2760), .Y(addr[24]) );
  TBUFX2TS \addr_calc/addr_tri4[20]  ( .A(\addr_calc/fir_write_addr[20] ), 
        .OE(n2761), .Y(addr[20]) );
  TBUFX2TS \addr_calc/addr_tri4[17]  ( .A(\addr_calc/fir_write_addr[17] ), 
        .OE(n2762), .Y(addr[17]) );
  TBUFX2TS \addr_calc/addr_tri4[14]  ( .A(\addr_calc/fir_write_addr[14] ), 
        .OE(n2763), .Y(addr[14]) );
  TBUFX2TS \addr_calc/addr_tri4[12]  ( .A(\addr_calc/fir_write_addr[12] ), 
        .OE(n2763), .Y(addr[12]) );
  TBUFX2TS \addr_calc/addr_tri4[11]  ( .A(\addr_calc/fir_write_addr[11] ), 
        .OE(n2764), .Y(addr[11]) );
  TBUFX2TS \addr_calc/addr_tri4[8]  ( .A(\addr_calc/fir_write_addr[8] ), .OE(
        n2764), .Y(addr[8]) );
  TBUFX2TS \addr_calc/addr_tri4[6]  ( .A(\addr_calc/fir_write_addr[6] ), .OE(
        n2765), .Y(addr[6]) );
  TBUFX2TS \addr_calc/addr_tri4[5]  ( .A(\addr_calc/fir_write_addr[5] ), .OE(
        n2765), .Y(addr[5]) );
  TBUFX2TS \addr_calc/addr_tri5[20]  ( .A(\addr_calc/iir_read_addr[20] ), .OE(
        n2769), .Y(addr[20]) );
  TBUFX2TS \addr_calc/addr_tri5[14]  ( .A(\addr_calc/iir_read_addr[14] ), .OE(
        n2771), .Y(addr[14]) );
  TBUFX2TS \addr_calc/addr_tri5[12]  ( .A(\addr_calc/iir_read_addr[12] ), .OE(
        n2771), .Y(addr[12]) );
  TBUFX2TS \addr_calc/addr_tri5[11]  ( .A(\addr_calc/iir_read_addr[11] ), .OE(
        n2772), .Y(addr[11]) );
  TBUFX2TS \addr_calc/addr_tri5[8]  ( .A(\addr_calc/iir_read_addr[8] ), .OE(
        n2772), .Y(addr[8]) );
  TBUFX2TS \addr_calc/addr_tri5[6]  ( .A(\addr_calc/iir_read_addr[6] ), .OE(
        n2773), .Y(addr[6]) );
  TBUFX2TS \addr_calc/addr_tri5[5]  ( .A(\addr_calc/iir_read_addr[5] ), .OE(
        n2773), .Y(addr[5]) );
  TBUFX2TS \addr_calc/addr_tri5[2]  ( .A(\addr_calc/iir_read_addr[2] ), .OE(
        n2774), .Y(addr[2]) );
  TBUFX2TS \addr_calc/addr_tri6[24]  ( .A(\addr_calc/iir_write_addr[24] ), 
        .OE(n2776), .Y(addr[24]) );
  TBUFX2TS \addr_calc/addr_tri6[20]  ( .A(\addr_calc/iir_write_addr[20] ), 
        .OE(n2777), .Y(addr[20]) );
  TBUFX2TS \addr_calc/addr_tri6[17]  ( .A(\addr_calc/iir_write_addr[17] ), 
        .OE(n2778), .Y(addr[17]) );
  TBUFX2TS \addr_calc/addr_tri6[14]  ( .A(\addr_calc/iir_write_addr[14] ), 
        .OE(n2779), .Y(addr[14]) );
  TBUFX2TS \addr_calc/addr_tri6[12]  ( .A(\addr_calc/iir_write_addr[12] ), 
        .OE(n2779), .Y(addr[12]) );
  TBUFX2TS \addr_calc/addr_tri6[11]  ( .A(\addr_calc/iir_write_addr[11] ), 
        .OE(n2780), .Y(addr[11]) );
  TBUFX2TS \addr_calc/addr_tri6[8]  ( .A(\addr_calc/iir_write_addr[8] ), .OE(
        n2780), .Y(addr[8]) );
  TBUFX2TS \addr_calc/addr_tri6[6]  ( .A(\addr_calc/iir_write_addr[6] ), .OE(
        n2781), .Y(addr[6]) );
  TBUFX2TS \addr_calc/addr_tri6[5]  ( .A(\addr_calc/iir_write_addr[5] ), .OE(
        n2781), .Y(addr[5]) );
  DFFQX2TS \addr_calc/fir_read_calc/counter/count_reg[28]  ( .D(n1070), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[28] ) );
  DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[2]  ( .D(n1128), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[2] ) );
  DFFQX1TS \addr_calc/fir_read_calc/counter/count_reg[29]  ( .D(n1069), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[29] ) );
  DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[0]  ( .D(n1098), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[0] ) );
  DFFHQX1TS \addr_calc/iir_read_calc/counter/count_reg[21]  ( .D(n950), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[21] ) );
  DFFHQX1TS \addr_calc/fir_write_calc/counter/count_reg[21]  ( .D(n1109), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[21] ) );
  DFFHQX1TS \addr_calc/fft_write_calc/counter/count_reg[21]  ( .D(n1045), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[21] ) );
  DFFHQX1TS \addr_calc/fft_read_calc/counter/count_reg[21]  ( .D(n1013), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[21] ) );
  DFFHQX1TS \addr_calc/fir_write_calc/counter/count_reg[15]  ( .D(n1115), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[15] ) );
  DFFHQX1TS \addr_calc/fir_write_calc/counter/count_reg[19]  ( .D(n1111), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[19] ) );
  DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[13]  ( .D(n1021), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[13] ) );
  DFFHQX1TS \addr_calc/fft_read_calc/counter/count_reg[17]  ( .D(n1017), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[17] ) );
  DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[10]  ( .D(n1088), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[10] ) );
  DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[16]  ( .D(n1082), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[16] ) );
  DFFQX1TS \pla_top/fir_enable_reg  ( .D(n1133), .CK(clk), .Q(n2814) );
  DFFHQX2TS \addr_calc/fft_write_calc/counter/count_reg[4]  ( .D(n1062), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[4] ) );
  DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[5]  ( .D(n966), .CK(clk), .Q(\addr_calc/iir_read_calc/count[5] ) );
  DFFQX2TS \addr_calc/iir_read_calc/counter/count_reg[30]  ( .D(n941), .CK(clk), .Q(\addr_calc/iir_read_calc/count[30] ) );
  DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[14]  ( .D(n1116), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[14] ) );
  DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[18]  ( .D(n1112), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[18] ) );
  DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[14]  ( .D(n1084), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[14] ) );
  DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[18]  ( .D(n1080), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[18] ) );
  DFFHQX2TS \addr_calc/fft_write_calc/counter/count_reg[18]  ( .D(n1048), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[18] ) );
  DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[14]  ( .D(n1020), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[14] ) );
  DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[18]  ( .D(n953), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[18] ) );
  DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[22]  ( .D(n1108), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[22] ) );
  DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[22]  ( .D(n1076), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[22] ) );
  DFFHQX2TS \addr_calc/fft_write_calc/counter/count_reg[22]  ( .D(n1044), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[22] ) );
  DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[22]  ( .D(n1012), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[22] ) );
  DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[20]  ( .D(n1110), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[20] ) );
  DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[20]  ( .D(n1078), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[20] ) );
  DFFHQX2TS \addr_calc/fft_write_calc/counter/count_reg[20]  ( .D(n1046), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[20] ) );
  DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[20]  ( .D(n951), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[20] ) );
  DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[12]  ( .D(n1022), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[12] ) );
  DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[0]  ( .D(n1034), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[0] ) );
  DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[7]  ( .D(n1027), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[7] ) );
  DFFHQX2TS \addr_calc/iir_write_calc/counter/count_reg[7]  ( .D(n995), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[7] ) );
  DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[9]  ( .D(n962), .CK(clk), .Q(\addr_calc/iir_read_calc/count[9] ) );
  DFFQX2TS \addr_calc/fir_read_calc/counter/count_reg[30]  ( .D(n1068), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[30] ) );
  DFFQX2TS \addr_calc/fft_write_calc/counter/count_reg[30]  ( .D(n1036), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[30] ) );
  DFFQX2TS \addr_calc/fft_read_calc/counter/count_reg[30]  ( .D(n1004), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[30] ) );
  TBUFX2TS \addr_calc/addr_tri[24]  ( .A(\addr_calc/fft_read_addr[24] ), .OE(
        n2736), .Y(addr[24]) );
  TBUFX2TS \addr_calc/addr_tri[20]  ( .A(\addr_calc/fft_read_addr[20] ), .OE(
        n2737), .Y(addr[20]) );
  TBUFX2TS \addr_calc/addr_tri[17]  ( .A(\addr_calc/fft_read_addr[17] ), .OE(
        n2738), .Y(addr[17]) );
  AOI21XLTS U346 ( .A0(fir_enable), .A1(n1828), .B0(n925), .Y(n924) );
  AOI32XLTS U23 ( .A0(fir_read_done), .A1(n2586), .A2(n2069), .B0(
        fft_read_done), .B1(fft_enable), .Y(n791) );
  AND2XLTS U342 ( .A(iir_put_req_reg), .B(n796), .Y(iir_put_req) );
  NOR3XLTS U351 ( .A(n2071), .B(n2061), .C(n900), .Y(n927) );
  OAI21XLTS U376 ( .A0(n2321), .A1(n2317), .B0(n2073), .Y(n939) );
  NOR2XLTS U358 ( .A(n2067), .B(n2071), .Y(\data_cntl/N266 ) );
  AOI21XLTS U362 ( .A0(iir_enable), .A1(n2061), .B0(fft_enable), .Y(
        \data_cntl/N263 ) );
  AOI21XLTS U383 ( .A0(n1861), .A1(n2060), .B0(n2072), .Y(n940) );
  AOI33XLTS U377 ( .A0(n2334), .A1(n2317), .A2(n2074), .B0(n2072), .B1(n2321), 
        .B2(n2319), .Y(\data_cntl/N250 ) );
  OAI21XLTS U359 ( .A0(n2063), .A1(fir_enable), .B0(n2586), .Y(
        \data_cntl/N260 ) );
  NOR3X1TS U352 ( .A(n1829), .B(n2060), .C(n925), .Y(n798) );
  NOR3X1TS U25 ( .A(n796), .B(n797), .C(n798), .Y(n790) );
  AOI31X1TS U21 ( .A0(n790), .A1(n791), .A2(n792), .B0(n793), .Y(
        ram_write_enable) );
  NOR2X1TS U314 ( .A(n2311), .B(n903), .Y(n872) );
  NOR2X1TS U311 ( .A(n2336), .B(n903), .Y(n902) );
  OAI21X1TS U303 ( .A0(fft_read_done), .A1(n1828), .B0(n887), .Y(n873) );
  AOI21X1TS U301 ( .A0(fir_write_done), .A1(n900), .B0(n884), .Y(n889) );
  AOI32X1TS U312 ( .A0(iir_write_done), .A1(n2055), .A2(n898), .B0(n899), .B1(
        n2054), .Y(n891) );
  NOR2X1TS U300 ( .A(n898), .B(n899), .Y(n893) );
  OAI31X1TS U298 ( .A0(n870), .A1(n895), .A2(n1828), .B0(n897), .Y(n894) );
  AOI32X1TS U297 ( .A0(n2054), .A1(n893), .A2(iir_write_done), .B0(n894), .B1(
        n2054), .Y(n892) );
  OAI31X1TS U296 ( .A0(n890), .A1(n889), .A2(n891), .B0(n892), .Y(n1134) );
  INVX2TS U307 ( .A(n2054), .Y(n869) );
  NOR3X1TS U295 ( .A(n887), .B(n888), .C(n889), .Y(n886) );
  OAI31X1TS U293 ( .A0(fir_write_done), .A1(n869), .A2(n884), .B0(n885), .Y(
        n1133) );
  OAI31X1TS U277 ( .A0(n1478), .A1(n869), .A2(n870), .B0(n871), .Y(n1131) );
  AND2XLTS U379 ( .A(\data_cntl/N265 ), .B(\data_cntl/N159 ), .Y(
        \addr_calc/N223 ) );
  AND2XLTS U387 ( .A(\data_cntl/N262 ), .B(\data_cntl/N95 ), .Y(
        \addr_calc/N219 ) );
  AND2XLTS U391 ( .A(\data_cntl/N259 ), .B(\data_cntl/N9 ), .Y(
        \addr_calc/N217 ) );
  NOR3X1TS U22 ( .A(\data_cntl/N267 ), .B(\data_cntl/N261 ), .C(
        \data_cntl/N264 ), .Y(n793) );
  NOR3X1TS U26 ( .A(\data_cntl/N262 ), .B(\data_cntl/N265 ), .C(
        \data_cntl/N259 ), .Y(n795) );
  NOR2X1TS U24 ( .A(n795), .B(n790), .Y(ram_read_enable) );
  NOR2BX1TS U327 ( .AN(chipselect), .B(n2116), .Y(n801) );
  AOI211XLTS U357 ( .A0(n1829), .A1(n895), .B0(n2587), .C0(n929), .Y(
        fft_get_req) );
  NOR4XLTS U325 ( .A(n2114), .B(n2095), .C(n2086), .D(n2105), .Y(n904) );
  NOR4XLTS U324 ( .A(n2110), .B(n2092), .C(n2084), .D(n2103), .Y(n905) );
  NOR4XLTS U339 ( .A(\addr_calc/iir_write_calc/count[23] ), .B(
        \addr_calc/iir_write_calc/count[22] ), .C(
        \addr_calc/iir_write_calc/count[21] ), .D(
        \addr_calc/iir_write_calc/count[20] ), .Y(n920) );
  NOR4XLTS U337 ( .A(n1951), .B(n1948), .C(n2570), .D(n1945), .Y(n922) );
  NOR4XLTS U72 ( .A(n2565), .B(\addr_calc/iir_read_calc/count[22] ), .C(n1687), 
        .D(\addr_calc/iir_read_calc/count[20] ), .Y(n815) );
  NOR4XLTS U151 ( .A(n1979), .B(\addr_calc/fft_read_calc/count[19] ), .C(
        \addr_calc/fft_read_calc/count[18] ), .D(n1960), .Y(n832) );
  NOR4XLTS U150 ( .A(\addr_calc/fft_read_calc/count[23] ), .B(n1665), .C(n1953), .D(\addr_calc/fft_read_calc/count[20] ), .Y(n833) );
  NOR4XLTS U275 ( .A(\addr_calc/fir_write_calc/count[23] ), .B(n1668), .C(
        n1892), .D(n1669), .Y(n866) );
  NOR4XLTS U273 ( .A(\addr_calc/fir_write_calc/count[16] ), .B(n1883), .C(
        \addr_calc/fir_write_calc/count[14] ), .D(
        \addr_calc/fir_write_calc/count[13] ), .Y(n868) );
  NOR4XLTS U290 ( .A(\addr_calc/fir_read_calc/count[23] ), .B(n1691), .C(n1879), .D(n1985), .Y(n881) );
  NOR4XLTS U340 ( .A(n1931), .B(\addr_calc/iir_write_calc/count[19] ), .C(
        n2571), .D(n1954), .Y(n919) );
  NOR4XLTS U73 ( .A(n1898), .B(n2556), .C(n2025), .D(
        \addr_calc/iir_read_calc/count[17] ), .Y(n814) );
  NOR4XLTS U196 ( .A(\addr_calc/fft_write_calc/count[23] ), .B(
        \addr_calc/fft_write_calc/count[22] ), .C(n1918), .D(
        \addr_calc/fft_write_calc/count[20] ), .Y(n847) );
  NOR4XLTS U276 ( .A(n1868), .B(\addr_calc/fir_write_calc/count[19] ), .C(
        n2006), .D(\addr_calc/fir_write_calc/count[17] ), .Y(n865) );
  INVX2TS U353 ( .A(n928), .Y(n925) );
  DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[25]  ( .D(n1041), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[25] ) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[17]  ( .D(n985), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[17] ) );
  DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[25]  ( .D(n1009), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[25] ) );
  TBUFX4TS \addr_calc/addr_tri3[30]  ( .A(\addr_calc/fir_read_addr[30] ), .OE(
        n2751), .Y(addr[30]) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[25]  ( .D(n977), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[25] ) );
  TBUFX12TS \addr_calc/addr_tri5[31]  ( .A(\addr_calc/iir_read_addr[31] ), 
        .OE(n2767), .Y(addr[31]) );
  DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[24]  ( .D(n1010), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[24] ) );
  DFFHQX8TS \addr_calc/fir_read_calc/counter/count_reg[25]  ( .D(n1073), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[25] ) );
  DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[24]  ( .D(n1042), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[24] ) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[16]  ( .D(n955), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[16] ) );
  TBUFX12TS \addr_calc/addr_tri3[31]  ( .A(\addr_calc/fir_read_addr[31] ), 
        .OE(n2751), .Y(addr[31]) );
  DFFHQX8TS \addr_calc/fir_read_calc/counter/count_reg[24]  ( .D(n1074), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[24] ) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[29]  ( .D(n942), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[29] ) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[19]  ( .D(n983), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[19] ) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[24]  ( .D(n947), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[24] ) );
  TBUFX4TS \addr_calc/addr_tri4[26]  ( .A(\addr_calc/fir_write_addr[26] ), 
        .OE(n2760), .Y(addr[26]) );
  TBUFX6TS \addr_calc/addr_tri4[30]  ( .A(\addr_calc/fir_write_addr[30] ), 
        .OE(n2759), .Y(addr[30]) );
  TBUFX12TS \addr_calc/addr_tri5[27]  ( .A(\addr_calc/iir_read_addr[27] ), 
        .OE(n2768), .Y(addr[27]) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[25]  ( .D(n946), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[25] ) );
  DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[29]  ( .D(n1037), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[29] ) );
  DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[29]  ( .D(n1005), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[29] ) );
  TBUFX6TS \addr_calc/addr_tri[21]  ( .A(\addr_calc/fft_read_addr[21] ), .OE(
        n2737), .Y(addr[21]) );
  TBUFX16TS \addr_calc/addr_tri4[31]  ( .A(\addr_calc/fir_write_addr[31] ), 
        .OE(n2759), .Y(addr[31]) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[0]  ( .D(n1002), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[0] ) );
  DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[3]  ( .D(n968), .CK(clk), .Q(\addr_calc/iir_read_calc/count[3] ) );
  TBUFX6TS \addr_calc/addr_tri[30]  ( .A(\addr_calc/fft_read_addr[30] ), .OE(
        n2735), .Y(addr[30]) );
  TBUFX4TS \addr_calc/addr_tri5[30]  ( .A(\addr_calc/iir_read_addr[30] ), .OE(
        n2767), .Y(addr[30]) );
  DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[0]  ( .D(n971), .CK(clk), .Q(\addr_calc/iir_read_calc/count[0] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[5]  ( .D(n997), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[5] ) );
  TBUFX16TS \addr_calc/addr_tri[31]  ( .A(\addr_calc/fft_read_addr[31] ), .OE(
        n2735), .Y(addr[31]) );
  DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[15]  ( .D(n1019), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[15] ) );
  TBUFX4TS \addr_calc/addr_tri6[15]  ( .A(\addr_calc/iir_write_addr[15] ), 
        .OE(n2779), .Y(addr[15]) );
  TBUFX4TS \addr_calc/addr_tri4[15]  ( .A(\addr_calc/fir_write_addr[15] ), 
        .OE(n2763), .Y(addr[15]) );
  DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[31]  ( .D(n1067), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[31] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[15]  ( .D(n1051), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[15] ) );
  DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[27]  ( .D(n1039), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[27] ) );
  TBUFX12TS \addr_calc/addr_tri4[23]  ( .A(\addr_calc/fir_write_addr[23] ), 
        .OE(n2761), .Y(addr[23]) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[19]  ( .D(n1015), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[19] ) );
  TBUFX4TS \addr_calc/addr_tri[26]  ( .A(\addr_calc/fft_read_addr[26] ), .OE(
        n2736), .Y(addr[26]) );
  TBUFX4TS \addr_calc/addr_tri5[26]  ( .A(\addr_calc/iir_read_addr[26] ), .OE(
        n2768), .Y(addr[26]) );
  TBUFX4TS \addr_calc/addr_tri6[26]  ( .A(\addr_calc/iir_write_addr[26] ), 
        .OE(n2776), .Y(addr[26]) );
  TBUFX4TS \addr_calc/addr_tri3[26]  ( .A(\addr_calc/fir_read_addr[26] ), .OE(
        n2752), .Y(addr[26]) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[9]  ( .D(n1121), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[9] ) );
  TBUFX4TS \addr_calc/addr_tri4[22]  ( .A(\addr_calc/fir_write_addr[22] ), 
        .OE(n2761), .Y(addr[22]) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[27]  ( .D(n975), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[27] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[29]  ( .D(n1101), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[29] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[6]  ( .D(n1060), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[6] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[13]  ( .D(n1053), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[13] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[21]  ( .D(n981), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[21] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[28]  ( .D(n974), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[28] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[27]  ( .D(n1103), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[27] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[17]  ( .D(n1113), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[17] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[5]  ( .D(n1125), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[5] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[11]  ( .D(n1055), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[11] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[27]  ( .D(n1007), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[27] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[19]  ( .D(n1047), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[19] ) );
  OAI21X1TS \add_x_19_4/U70  ( .A0(\add_x_19_4/n78 ), .A1(\add_x_19_4/n82 ), 
        .B0(\add_x_19_4/n79 ), .Y(\add_x_19_4/n77 ) );
  NAND2X1TS \add_x_19_4/U255  ( .A(\addr_calc/iir_read_calc/count[0] ), .B(
        n2392), .Y(\add_x_19_4/n191 ) );
  XOR2X1TS \add_x_19_4/U244  ( .A(\add_x_19_4/n31 ), .B(\add_x_19_4/n191 ), 
        .Y(\addr_calc/iir_read_addr[1] ) );
  XOR2X1TS \add_x_19_4/U238  ( .A(\add_x_19_4/n186 ), .B(\add_x_19_4/n30 ), 
        .Y(\addr_calc/iir_read_addr[2] ) );
  AOI21X1TS \add_x_19_4/U214  ( .A0(\add_x_19_4/n177 ), .A1(\add_x_19_4/n168 ), 
        .B0(\add_x_19_4/n169 ), .Y(\add_x_19_4/n167 ) );
  AOI21X1TS \add_x_19_4/U173  ( .A0(\add_x_19_4/n146 ), .A1(\add_x_19_4/n213 ), 
        .B0(\add_x_19_4/n143 ), .Y(\add_x_19_4/n141 ) );
  OAI21X1TS \add_x_19_4/U181  ( .A0(\add_x_19_4/n156 ), .A1(\add_x_19_4/n147 ), 
        .B0(\add_x_19_4/n148 ), .Y(\add_x_19_4/n146 ) );
  OAI21X1TS \add_x_19_4/U156  ( .A0(\add_x_19_4/n133 ), .A1(\add_x_19_4/n131 ), 
        .B0(\add_x_19_4/n132 ), .Y(\add_x_19_4/n130 ) );
  AOI21X1TS \add_x_19_4/U121  ( .A0(\add_x_19_4/n112 ), .A1(\add_x_19_4/n207 ), 
        .B0(\add_x_19_4/n109 ), .Y(\add_x_19_4/n107 ) );
  OAI21X1TS \add_x_19_4/U90  ( .A0(\add_x_19_4/n91 ), .A1(\add_x_19_4/n89 ), 
        .B0(\add_x_19_4/n90 ), .Y(\add_x_19_4/n88 ) );
  NOR2X1TS \add_x_19_4/U10  ( .A(n1684), .B(n2456), .Y(\add_x_19_4/n36 ) );
  AOI21X1TS \add_x_19_4/U33  ( .A0(\add_x_19_4/n53 ), .A1(\add_x_19_4/n62 ), 
        .B0(\add_x_19_4/n54 ), .Y(\add_x_19_4/n52 ) );
  OAI21X1TS \add_x_19_4/U35  ( .A0(\add_x_19_4/n55 ), .A1(\add_x_19_4/n59 ), 
        .B0(\add_x_19_4/n56 ), .Y(\add_x_19_4/n54 ) );
  OAI21X1TS \add_x_19_4/U49  ( .A0(\add_x_19_4/n63 ), .A1(\add_x_19_4/n67 ), 
        .B0(\add_x_19_4/n64 ), .Y(\add_x_19_4/n62 ) );
  OAI21X1TS \add_x_19_4/U84  ( .A0(\add_x_19_4/n86 ), .A1(\add_x_19_4/n90 ), 
        .B0(\add_x_19_4/n87 ), .Y(\add_x_19_4/n85 ) );
  AOI21X1TS \add_x_19_4/U99  ( .A0(\add_x_19_4/n95 ), .A1(\add_x_19_4/n104 ), 
        .B0(\add_x_19_4/n96 ), .Y(\add_x_19_4/n94 ) );
  OAI21X1TS \add_x_19_4/U101  ( .A0(\add_x_19_4/n97 ), .A1(\add_x_19_4/n101 ), 
        .B0(\add_x_19_4/n98 ), .Y(\add_x_19_4/n96 ) );
  OAI21X1TS \add_x_19_4/U115  ( .A0(\add_x_19_4/n105 ), .A1(\add_x_19_4/n111 ), 
        .B0(\add_x_19_4/n106 ), .Y(\add_x_19_4/n104 ) );
  NOR2X1TS \add_x_19_4/U24  ( .A(\add_x_19_4/n51 ), .B(\add_x_19_4/n48 ), .Y(
        \add_x_19_4/n46 ) );
  NOR2X1TS \add_x_19_4/U34  ( .A(\add_x_19_4/n58 ), .B(\add_x_19_4/n55 ), .Y(
        \add_x_19_4/n53 ) );
  NOR2X1TS \add_x_19_4/U83  ( .A(\add_x_19_4/n89 ), .B(\add_x_19_4/n86 ), .Y(
        \add_x_19_4/n84 ) );
  NOR2X1TS \add_x_19_4/U100  ( .A(\add_x_19_4/n100 ), .B(\add_x_19_4/n97 ), 
        .Y(\add_x_19_4/n95 ) );
  NOR2X1TS \add_x_19_4/U114  ( .A(\add_x_19_4/n110 ), .B(\add_x_19_4/n105 ), 
        .Y(\add_x_19_4/n103 ) );
  OAI21X1TS \add_x_19_4/U167  ( .A0(\add_x_19_4/n139 ), .A1(\add_x_19_4/n145 ), 
        .B0(\add_x_19_4/n140 ), .Y(\add_x_19_4/n138 ) );
  OAI21X1TS \add_x_19_4/U185  ( .A0(\add_x_19_4/n151 ), .A1(\add_x_19_4/n155 ), 
        .B0(\add_x_19_4/n152 ), .Y(\add_x_19_4/n150 ) );
  NOR2X1TS \add_x_19_4/U166  ( .A(\add_x_19_4/n144 ), .B(\add_x_19_4/n139 ), 
        .Y(\add_x_19_4/n137 ) );
  NOR2X1TS \add_x_19_4/U184  ( .A(\add_x_19_4/n154 ), .B(\add_x_19_4/n151 ), 
        .Y(\add_x_19_4/n149 ) );
  NOR2X1TS \add_x_19_4/U201  ( .A(\add_x_19_4/n165 ), .B(\add_x_19_4/n162 ), 
        .Y(\add_x_19_4/n160 ) );
  NOR2X1TS \add_x_19_4/U215  ( .A(\add_x_19_4/n175 ), .B(\add_x_19_4/n170 ), 
        .Y(\add_x_19_4/n168 ) );
  NOR2X1TS \add_x_19_4/U249  ( .A(\addr_calc/iir_read_calc/count[1] ), .B(
        n2453), .Y(\add_x_19_4/n188 ) );
  XOR2X1TS \add_x_19_4/U207  ( .A(\add_x_19_4/n167 ), .B(\add_x_19_4/n26 ), 
        .Y(\addr_calc/iir_read_addr[6] ) );
  XOR2X1TS \add_x_19_4/U161  ( .A(\add_x_19_4/n141 ), .B(\add_x_19_4/n21 ), 
        .Y(\addr_calc/iir_read_addr[11] ) );
  XOR2X1TS \add_x_19_4/U112  ( .A(\add_x_19_4/n107 ), .B(\add_x_19_4/n15 ), 
        .Y(\addr_calc/iir_read_addr[17] ) );
  NAND2X1TS \add_x_19_4/U11  ( .A(n1684), .B(n2458), .Y(\add_x_19_4/n37 ) );
  NAND2X1TS \add_x_19_4/U19  ( .A(n1840), .B(n2388), .Y(\add_x_19_4/n42 ) );
  NAND2X1TS \add_x_19_4/U29  ( .A(n2561), .B(n2384), .Y(\add_x_19_4/n49 ) );
  NAND2X1TS \add_x_19_4/U39  ( .A(n1929), .B(n2498), .Y(\add_x_19_4/n56 ) );
  NAND2X1TS \add_x_19_4/U45  ( .A(\addr_calc/iir_read_calc/count[26] ), .B(
        n2378), .Y(\add_x_19_4/n59 ) );
  NAND2X1TS \add_x_19_4/U53  ( .A(n1926), .B(n2491), .Y(\add_x_19_4/n64 ) );
  NAND2X1TS \add_x_19_4/U59  ( .A(n2034), .B(n2462), .Y(\add_x_19_4/n67 ) );
  NAND2X1TS \add_x_19_4/U74  ( .A(\addr_calc/iir_read_calc/count[23] ), .B(
        n2470), .Y(\add_x_19_4/n79 ) );
  NAND2X1TS \add_x_19_4/U80  ( .A(\addr_calc/iir_read_calc/count[22] ), .B(
        n2465), .Y(\add_x_19_4/n82 ) );
  NAND2X1TS \add_x_19_4/U88  ( .A(n1687), .B(n2449), .Y(\add_x_19_4/n87 ) );
  NAND2X1TS \add_x_19_4/U94  ( .A(n2028), .B(n2442), .Y(\add_x_19_4/n90 ) );
  NAND2X1TS \add_x_19_4/U105  ( .A(\addr_calc/iir_read_calc/count[19] ), .B(
        n2489), .Y(\add_x_19_4/n98 ) );
  NAND2X1TS \add_x_19_4/U111  ( .A(n2025), .B(n2434), .Y(\add_x_19_4/n101 ) );
  NAND2X1TS \add_x_19_4/U127  ( .A(n1916), .B(n2401), .Y(\add_x_19_4/n111 ) );
  NOR2X1TS \add_x_19_4/U58  ( .A(\addr_calc/iir_read_calc/count[24] ), .B(
        n2460), .Y(\add_x_19_4/n66 ) );
  NOR2X1TS \add_x_19_4/U87  ( .A(n1687), .B(n2448), .Y(\add_x_19_4/n86 ) );
  NOR2X1TS \add_x_19_4/U93  ( .A(n2028), .B(n2440), .Y(\add_x_19_4/n89 ) );
  NOR2X1TS \add_x_19_4/U110  ( .A(n2025), .B(n2434), .Y(\add_x_19_4/n100 ) );
  NOR2X1TS \add_x_19_4/U118  ( .A(n1920), .B(n2481), .Y(\add_x_19_4/n105 ) );
  NOR2X1TS \add_x_19_4/U126  ( .A(n1916), .B(n2400), .Y(\add_x_19_4/n110 ) );
  NAND2X1TS \add_x_19_4/U140  ( .A(\addr_calc/iir_read_calc/count[15] ), .B(
        n2477), .Y(\add_x_19_4/n121 ) );
  NAND2X1TS \add_x_19_4/U154  ( .A(\addr_calc/iir_read_calc/count[13] ), .B(
        n2416), .Y(\add_x_19_4/n129 ) );
  NAND2X1TS \add_x_19_4/U179  ( .A(n1909), .B(n2412), .Y(\add_x_19_4/n145 ) );
  NAND2X1TS \add_x_19_4/U189  ( .A(n1685), .B(n1980), .Y(\add_x_19_4/n152 ) );
  NAND2X1TS \add_x_19_4/U195  ( .A(\addr_calc/iir_read_calc/count[8] ), .B(
        n1864), .Y(\add_x_19_4/n155 ) );
  NOR2X1TS \add_x_19_4/U153  ( .A(\addr_calc/iir_read_calc/count[13] ), .B(
        n2416), .Y(\add_x_19_4/n128 ) );
  NOR2X1TS \add_x_19_4/U178  ( .A(n1909), .B(n2412), .Y(\add_x_19_4/n144 ) );
  NOR2X1TS \add_x_19_4/U194  ( .A(\addr_calc/iir_read_calc/count[8] ), .B(
        n1864), .Y(\add_x_19_4/n154 ) );
  NAND2X1TS \add_x_19_4/U206  ( .A(n1905), .B(n2420), .Y(\add_x_19_4/n163 ) );
  NAND2X1TS \add_x_19_4/U212  ( .A(n2428), .B(
        \addr_calc/iir_read_calc/count[6] ), .Y(\add_x_19_4/n166 ) );
  NAND2X1TS \add_x_19_4/U228  ( .A(\addr_calc/iir_read_calc/count[4] ), .B(
        n2398), .Y(\add_x_19_4/n176 ) );
  NOR2X1TS \add_x_19_4/U211  ( .A(\addr_calc/iir_read_calc/count[6] ), .B(
        n2430), .Y(\add_x_19_4/n165 ) );
  NOR2X1TS \add_x_19_4/U227  ( .A(\addr_calc/iir_read_calc/count[4] ), .B(
        n2398), .Y(\add_x_19_4/n175 ) );
  NAND2X1TS \add_x_19_4/U237  ( .A(n1902), .B(n2438), .Y(\add_x_19_4/n182 ) );
  NAND2X1TS \add_x_19_4/U250  ( .A(\addr_calc/iir_read_calc/count[1] ), .B(
        n2454), .Y(\add_x_19_4/n189 ) );
  NOR2X1TS \add_x_19_4/U242  ( .A(\addr_calc/iir_read_calc/count[2] ), .B(
        n2445), .Y(\add_x_19_4/n184 ) );
  NAND2X1TS \add_x_19_4/U247  ( .A(\add_x_19_4/n222 ), .B(\add_x_19_4/n189 ), 
        .Y(\add_x_19_4/n31 ) );
  NAND2X1TS \add_x_19_4/U240  ( .A(\add_x_19_4/n221 ), .B(\add_x_19_4/n185 ), 
        .Y(\add_x_19_4/n30 ) );
  XNOR2X1TS \add_x_19_4/U221  ( .A(\add_x_19_4/n177 ), .B(\add_x_19_4/n28 ), 
        .Y(\addr_calc/iir_read_addr[4] ) );
  NAND2X1TS \add_x_19_4/U225  ( .A(\add_x_19_4/n219 ), .B(\add_x_19_4/n176 ), 
        .Y(\add_x_19_4/n28 ) );
  NAND2X1TS \add_x_19_4/U209  ( .A(\add_x_19_4/n217 ), .B(\add_x_19_4/n166 ), 
        .Y(\add_x_19_4/n26 ) );
  XNOR2X1TS \add_x_19_4/U172  ( .A(\add_x_19_4/n146 ), .B(\add_x_19_4/n22 ), 
        .Y(\addr_calc/iir_read_addr[10] ) );
  NAND2X1TS \add_x_19_4/U176  ( .A(\add_x_19_4/n213 ), .B(\add_x_19_4/n145 ), 
        .Y(\add_x_19_4/n22 ) );
  NAND2X1TS \add_x_19_4/U168  ( .A(\add_x_19_4/n212 ), .B(\add_x_19_4/n140 ), 
        .Y(\add_x_19_4/n21 ) );
  XNOR2X1TS \add_x_19_4/U147  ( .A(\add_x_19_4/n130 ), .B(\add_x_19_4/n19 ), 
        .Y(\addr_calc/iir_read_addr[13] ) );
  NAND2X1TS \add_x_19_4/U151  ( .A(n1632), .B(\add_x_19_4/n129 ), .Y(
        \add_x_19_4/n19 ) );
  NAND2X1TS \add_x_19_4/U116  ( .A(\add_x_19_4/n206 ), .B(\add_x_19_4/n106 ), 
        .Y(\add_x_19_4/n15 ) );
  XNOR2X1TS \add_x_19_4/U12  ( .A(\add_x_19_4/n43 ), .B(\add_x_19_4/n3 ), .Y(
        \addr_calc/iir_read_addr[29] ) );
  NAND2X1TS \add_x_19_4/U16  ( .A(n2634), .B(\add_x_19_4/n42 ), .Y(
        \add_x_19_4/n3 ) );
  NAND2X1TS \add_x_19_4/U102  ( .A(\add_x_19_4/n204 ), .B(\add_x_19_4/n98 ), 
        .Y(\add_x_19_4/n13 ) );
  NAND2X1TS \add_x_19_4/U85  ( .A(\add_x_19_4/n202 ), .B(\add_x_19_4/n87 ), 
        .Y(\add_x_19_4/n11 ) );
  NAND2X1TS \add_x_19_4/U36  ( .A(\add_x_19_4/n196 ), .B(\add_x_19_4/n56 ), 
        .Y(\add_x_19_4/n5 ) );
  NAND2X1TS \add_x_19_4/U119  ( .A(n1920), .B(n2480), .Y(\add_x_19_4/n106 ) );
  NAND2X1TS \add_x_19_4/U32  ( .A(\add_x_19_4/n61 ), .B(\add_x_19_4/n53 ), .Y(
        \add_x_19_4/n51 ) );
  NAND2X1TS \add_x_19_4/U98  ( .A(\add_x_19_4/n103 ), .B(\add_x_19_4/n95 ), 
        .Y(\add_x_19_4/n93 ) );
  NAND2X1TS \add_x_19_4/U171  ( .A(n1911), .B(n2406), .Y(\add_x_19_4/n140 ) );
  NAND2X1TS \add_x_19_4/U164  ( .A(\add_x_19_4/n149 ), .B(\add_x_19_4/n137 ), 
        .Y(\add_x_19_4/n135 ) );
  NAND2X1TS \add_x_19_4/U220  ( .A(\addr_calc/iir_read_calc/count[5] ), .B(
        n2483), .Y(\add_x_19_4/n171 ) );
  NOR2X1TS \add_x_19_2/U236  ( .A(\addr_calc/fir_read_calc/count[3] ), .B(
        n2437), .Y(\add_x_19_2/n181 ) );
  NOR2X1TS \add_x_19_2/U211  ( .A(\addr_calc/fir_read_calc/count[6] ), .B(
        n2430), .Y(\add_x_19_2/n165 ) );
  OAI21X1TS \add_x_19_2/U35  ( .A0(\add_x_19_2/n55 ), .A1(\add_x_19_2/n59 ), 
        .B0(\add_x_19_2/n56 ), .Y(\add_x_19_2/n54 ) );
  NAND2X1TS \add_x_19_2/U255  ( .A(\addr_calc/fir_read_calc/count[0] ), .B(
        n2392), .Y(\add_x_19_2/n191 ) );
  OAI21X1TS \add_x_19_2/U208  ( .A0(\add_x_19_2/n167 ), .A1(\add_x_19_2/n165 ), 
        .B0(\add_x_19_2/n166 ), .Y(\add_x_19_2/n164 ) );
  AOI21X1TS \add_x_19_2/U214  ( .A0(\add_x_19_2/n177 ), .A1(\add_x_19_2/n168 ), 
        .B0(\add_x_19_2/n169 ), .Y(\add_x_19_2/n167 ) );
  OAI21X1TS \add_x_19_2/U181  ( .A0(\add_x_19_2/n156 ), .A1(\add_x_19_2/n147 ), 
        .B0(\add_x_19_2/n148 ), .Y(\add_x_19_2/n146 ) );
  OAI21X1TS \add_x_19_2/U156  ( .A0(\add_x_19_2/n133 ), .A1(\add_x_19_2/n131 ), 
        .B0(\add_x_19_2/n132 ), .Y(\add_x_19_2/n130 ) );
  AOI21X1TS \add_x_19_2/U121  ( .A0(\add_x_19_2/n112 ), .A1(\add_x_19_2/n207 ), 
        .B0(\add_x_19_2/n109 ), .Y(\add_x_19_2/n107 ) );
  OAI21X1TS \add_x_19_2/U142  ( .A0(\add_x_19_2/n125 ), .A1(\add_x_19_2/n123 ), 
        .B0(\add_x_19_2/n124 ), .Y(\add_x_19_2/n122 ) );
  AOI21X1TS \add_x_19_2/U148  ( .A0(\add_x_19_2/n134 ), .A1(\add_x_19_2/n126 ), 
        .B0(\add_x_19_2/n127 ), .Y(\add_x_19_2/n125 ) );
  OAI21X1TS \add_x_19_2/U107  ( .A0(\add_x_19_2/n102 ), .A1(\add_x_19_2/n100 ), 
        .B0(\add_x_19_2/n101 ), .Y(\add_x_19_2/n99 ) );
  AOI21X1TS \add_x_19_2/U113  ( .A0(\add_x_19_2/n112 ), .A1(\add_x_19_2/n103 ), 
        .B0(\add_x_19_2/n104 ), .Y(\add_x_19_2/n102 ) );
  NOR2X1TS \add_x_19_2/U10  ( .A(n1838), .B(n2457), .Y(\add_x_19_2/n36 ) );
  AOI21X1TS \add_x_19_2/U33  ( .A0(\add_x_19_2/n53 ), .A1(\add_x_19_2/n62 ), 
        .B0(\add_x_19_2/n54 ), .Y(\add_x_19_2/n52 ) );
  OAI21X1TS \add_x_19_2/U49  ( .A0(\add_x_19_2/n63 ), .A1(\add_x_19_2/n67 ), 
        .B0(\add_x_19_2/n64 ), .Y(\add_x_19_2/n62 ) );
  AOI21X1TS \add_x_19_2/U99  ( .A0(\add_x_19_2/n95 ), .A1(\add_x_19_2/n104 ), 
        .B0(\add_x_19_2/n96 ), .Y(\add_x_19_2/n94 ) );
  OAI21X1TS \add_x_19_2/U101  ( .A0(\add_x_19_2/n97 ), .A1(\add_x_19_2/n101 ), 
        .B0(\add_x_19_2/n98 ), .Y(\add_x_19_2/n96 ) );
  OAI21X1TS \add_x_19_2/U115  ( .A0(\add_x_19_2/n105 ), .A1(\add_x_19_2/n111 ), 
        .B0(\add_x_19_2/n106 ), .Y(\add_x_19_2/n104 ) );
  NOR2X1TS \add_x_19_2/U48  ( .A(\add_x_19_2/n66 ), .B(\add_x_19_2/n63 ), .Y(
        \add_x_19_2/n61 ) );
  NOR2X1TS \add_x_19_2/U58  ( .A(n1983), .B(n2461), .Y(\add_x_19_2/n66 ) );
  NOR2X1TS \add_x_19_2/U65  ( .A(\add_x_19_2/n93 ), .B(\add_x_19_2/n74 ), .Y(
        \add_x_19_2/n72 ) );
  NOR2X1TS \add_x_19_2/U83  ( .A(\add_x_19_2/n89 ), .B(\add_x_19_2/n86 ), .Y(
        \add_x_19_2/n84 ) );
  NOR2X1TS \add_x_19_2/U100  ( .A(\add_x_19_2/n100 ), .B(\add_x_19_2/n97 ), 
        .Y(\add_x_19_2/n95 ) );
  NOR2X1TS \add_x_19_2/U114  ( .A(\add_x_19_2/n110 ), .B(\add_x_19_2/n105 ), 
        .Y(\add_x_19_2/n103 ) );
  OAI21X1TS \add_x_19_2/U150  ( .A0(\add_x_19_2/n128 ), .A1(\add_x_19_2/n132 ), 
        .B0(\add_x_19_2/n129 ), .Y(\add_x_19_2/n127 ) );
  NOR2X1TS \add_x_19_2/U139  ( .A(\addr_calc/fir_read_calc/count[15] ), .B(
        n2475), .Y(\add_x_19_2/n120 ) );
  NOR2X1TS \add_x_19_2/U149  ( .A(\add_x_19_2/n131 ), .B(\add_x_19_2/n128 ), 
        .Y(\add_x_19_2/n126 ) );
  NOR2X1TS \add_x_19_2/U166  ( .A(\add_x_19_2/n144 ), .B(\add_x_19_2/n139 ), 
        .Y(\add_x_19_2/n137 ) );
  NOR2X1TS \add_x_19_2/U170  ( .A(\addr_calc/fir_read_calc/count[11] ), .B(
        n2404), .Y(\add_x_19_2/n139 ) );
  NOR2X1TS \add_x_19_2/U184  ( .A(\add_x_19_2/n154 ), .B(\add_x_19_2/n151 ), 
        .Y(\add_x_19_2/n149 ) );
  NOR2X1TS \add_x_19_2/U215  ( .A(\add_x_19_2/n175 ), .B(\add_x_19_2/n170 ), 
        .Y(\add_x_19_2/n168 ) );
  OAI21X1TS \add_x_19_2/U246  ( .A0(\add_x_19_2/n188 ), .A1(\add_x_19_2/n191 ), 
        .B0(\add_x_19_2/n189 ), .Y(\add_x_19_2/n187 ) );
  NOR2X1TS \add_x_19_2/U249  ( .A(n1910), .B(n2453), .Y(\add_x_19_2/n188 ) );
  XOR2X1TS \add_x_19_2/U112  ( .A(\add_x_19_2/n107 ), .B(\add_x_19_2/n15 ), 
        .Y(\addr_calc/fir_read_addr[17] ) );
  NAND2X1TS \add_x_19_2/U11  ( .A(\addr_calc/fir_read_calc/count[30] ), .B(
        n2458), .Y(\add_x_19_2/n37 ) );
  NAND2X1TS \add_x_19_2/U19  ( .A(n1842), .B(n2390), .Y(\add_x_19_2/n42 ) );
  NAND2X1TS \add_x_19_2/U29  ( .A(n1871), .B(n2385), .Y(\add_x_19_2/n49 ) );
  NAND2X1TS \add_x_19_2/U39  ( .A(\addr_calc/fir_read_calc/count[27] ), .B(
        n2499), .Y(\add_x_19_2/n56 ) );
  NAND2X1TS \add_x_19_2/U45  ( .A(\addr_calc/fir_read_calc/count[26] ), .B(
        n2377), .Y(\add_x_19_2/n59 ) );
  NAND2X1TS \add_x_19_2/U53  ( .A(n1876), .B(n2493), .Y(\add_x_19_2/n64 ) );
  NAND2X1TS \add_x_19_2/U59  ( .A(n1983), .B(n2460), .Y(\add_x_19_2/n67 ) );
  NAND2X1TS \add_x_19_2/U74  ( .A(\addr_calc/fir_read_calc/count[23] ), .B(
        n2470), .Y(\add_x_19_2/n79 ) );
  NAND2X1TS \add_x_19_2/U80  ( .A(\addr_calc/fir_read_calc/count[22] ), .B(
        n2466), .Y(\add_x_19_2/n82 ) );
  NAND2X1TS \add_x_19_2/U88  ( .A(n1879), .B(n2448), .Y(\add_x_19_2/n87 ) );
  NAND2X1TS \add_x_19_2/U94  ( .A(n1985), .B(n2441), .Y(\add_x_19_2/n90 ) );
  NAND2X1TS \add_x_19_2/U105  ( .A(\addr_calc/fir_read_calc/count[19] ), .B(
        n2488), .Y(\add_x_19_2/n98 ) );
  NAND2X1TS \add_x_19_2/U111  ( .A(n1988), .B(n2433), .Y(\add_x_19_2/n101 ) );
  NAND2X1TS \add_x_19_2/U127  ( .A(n1888), .B(n2400), .Y(\add_x_19_2/n111 ) );
  NOR2X1TS \add_x_19_2/U52  ( .A(n1876), .B(n2491), .Y(\add_x_19_2/n63 ) );
  NOR2X1TS \add_x_19_2/U79  ( .A(n1691), .B(n2464), .Y(\add_x_19_2/n81 ) );
  NOR2X1TS \add_x_19_2/U93  ( .A(n1985), .B(n2442), .Y(\add_x_19_2/n89 ) );
  NOR2X1TS \add_x_19_2/U104  ( .A(\addr_calc/fir_read_calc/count[19] ), .B(
        n2487), .Y(\add_x_19_2/n97 ) );
  NOR2X1TS \add_x_19_2/U110  ( .A(n1988), .B(n2432), .Y(\add_x_19_2/n100 ) );
  NOR2X1TS \add_x_19_2/U118  ( .A(\addr_calc/fir_read_calc/count[17] ), .B(
        n2479), .Y(\add_x_19_2/n105 ) );
  NOR2X1TS \add_x_19_2/U126  ( .A(n1888), .B(n2401), .Y(\add_x_19_2/n110 ) );
  NAND2X1TS \add_x_19_2/U140  ( .A(\addr_calc/fir_read_calc/count[15] ), .B(
        n2476), .Y(\add_x_19_2/n121 ) );
  NAND2X1TS \add_x_19_2/U146  ( .A(\addr_calc/fir_read_calc/count[14] ), .B(
        n2424), .Y(\add_x_19_2/n124 ) );
  NAND2X1TS \add_x_19_2/U154  ( .A(\addr_calc/fir_read_calc/count[13] ), .B(
        n2417), .Y(\add_x_19_2/n129 ) );
  NAND2X1TS \add_x_19_2/U160  ( .A(\addr_calc/fir_read_calc/count[12] ), .B(
        n2409), .Y(\add_x_19_2/n132 ) );
  NAND2X1TS \add_x_19_2/U189  ( .A(n1900), .B(n2496), .Y(\add_x_19_2/n152 ) );
  NAND2X1TS \add_x_19_2/U195  ( .A(\addr_calc/fir_read_calc/count[8] ), .B(
        n2473), .Y(\add_x_19_2/n155 ) );
  NOR2X1TS \add_x_19_2/U153  ( .A(\addr_calc/fir_read_calc/count[13] ), .B(
        n2416), .Y(\add_x_19_2/n128 ) );
  NOR2X1TS \add_x_19_2/U159  ( .A(\addr_calc/fir_read_calc/count[12] ), .B(
        n2408), .Y(\add_x_19_2/n131 ) );
  NOR2X1TS \add_x_19_2/U194  ( .A(\addr_calc/fir_read_calc/count[8] ), .B(
        n2472), .Y(\add_x_19_2/n154 ) );
  NAND2X1TS \add_x_19_2/U212  ( .A(\addr_calc/fir_read_calc/count[6] ), .B(
        n2429), .Y(\add_x_19_2/n166 ) );
  NAND2X1TS \add_x_19_2/U228  ( .A(\addr_calc/fir_read_calc/count[4] ), .B(
        n2398), .Y(\add_x_19_2/n176 ) );
  NAND2X1TS \add_x_19_2/U237  ( .A(\addr_calc/fir_read_calc/count[3] ), .B(
        n2438), .Y(\add_x_19_2/n182 ) );
  NAND2X1TS \add_x_19_2/U243  ( .A(\addr_calc/fir_read_calc/count[2] ), .B(
        n2446), .Y(\add_x_19_2/n185 ) );
  NAND2X1TS \add_x_19_2/U250  ( .A(n1910), .B(n2452), .Y(\add_x_19_2/n189 ) );
  NOR2X1TS \add_x_19_2/U242  ( .A(\addr_calc/fir_read_calc/count[2] ), .B(
        n2446), .Y(\add_x_19_2/n184 ) );
  XNOR2X1TS \add_x_19_2/U221  ( .A(\add_x_19_2/n177 ), .B(\add_x_19_2/n28 ), 
        .Y(\addr_calc/fir_read_addr[4] ) );
  NAND2X1TS \add_x_19_2/U225  ( .A(\add_x_19_2/n219 ), .B(\add_x_19_2/n176 ), 
        .Y(\add_x_19_2/n28 ) );
  XNOR2X1TS \add_x_19_2/U196  ( .A(\add_x_19_2/n164 ), .B(\add_x_19_2/n25 ), 
        .Y(\addr_calc/fir_read_addr[7] ) );
  NAND2X1TS \add_x_19_2/U203  ( .A(\add_x_19_2/n216 ), .B(\add_x_19_2/n163 ), 
        .Y(\add_x_19_2/n25 ) );
  NAND2X1TS \add_x_19_2/U192  ( .A(\add_x_19_2/n215 ), .B(\add_x_19_2/n155 ), 
        .Y(\add_x_19_2/n24 ) );
  XNOR2X1TS \add_x_19_2/U147  ( .A(\add_x_19_2/n130 ), .B(\add_x_19_2/n19 ), 
        .Y(\addr_calc/fir_read_addr[13] ) );
  NAND2X1TS \add_x_19_2/U151  ( .A(\add_x_19_2/n210 ), .B(\add_x_19_2/n129 ), 
        .Y(\add_x_19_2/n19 ) );
  NAND2X1TS \add_x_19_2/U116  ( .A(\add_x_19_2/n206 ), .B(\add_x_19_2/n106 ), 
        .Y(\add_x_19_2/n15 ) );
  NAND2X1TS \add_x_19_2/U137  ( .A(\add_x_19_2/n208 ), .B(\add_x_19_2/n121 ), 
        .Y(\add_x_19_2/n17 ) );
  NAND2X1TS \add_x_19_2/U119  ( .A(\addr_calc/fir_read_calc/count[17] ), .B(
        n2479), .Y(\add_x_19_2/n106 ) );
  NAND2X1TS \add_x_19_2/U32  ( .A(\add_x_19_2/n61 ), .B(\add_x_19_2/n53 ), .Y(
        \add_x_19_2/n51 ) );
  NAND2X1TS \add_x_19_2/U98  ( .A(\add_x_19_2/n103 ), .B(\add_x_19_2/n95 ), 
        .Y(\add_x_19_2/n93 ) );
  NAND2X1TS \add_x_19_2/U171  ( .A(\addr_calc/fir_read_calc/count[11] ), .B(
        n2405), .Y(\add_x_19_2/n140 ) );
  NAND2X1TS \add_x_19_2/U133  ( .A(\add_x_19_2/n126 ), .B(\add_x_19_2/n118 ), 
        .Y(\add_x_19_2/n116 ) );
  NAND2X1TS \add_x_19_2/U164  ( .A(\add_x_19_2/n149 ), .B(\add_x_19_2/n137 ), 
        .Y(\add_x_19_2/n135 ) );
  NAND2X1TS \add_x_19_2/U220  ( .A(n1904), .B(n2484), .Y(\add_x_19_2/n171 ) );
  NOR2X1TS \add_x_19_1/U236  ( .A(\addr_calc/fft_write_calc/count[3] ), .B(
        n2436), .Y(\add_x_19_1/n181 ) );
  NOR2X1TS \add_x_19_1/U205  ( .A(\addr_calc/fft_write_calc/count[7] ), .B(
        n2421), .Y(\add_x_19_1/n162 ) );
  OAI21X1TS \add_x_19_1/U70  ( .A0(\add_x_19_1/n78 ), .A1(\add_x_19_1/n82 ), 
        .B0(\add_x_19_1/n79 ), .Y(\add_x_19_1/n77 ) );
  NAND2X1TS \add_x_19_1/U255  ( .A(n2035), .B(n2392), .Y(\add_x_19_1/n191 ) );
  AOI21X1TS \add_x_19_1/U222  ( .A0(\add_x_19_1/n177 ), .A1(\add_x_19_1/n219 ), 
        .B0(\add_x_19_1/n174 ), .Y(\add_x_19_1/n172 ) );
  AOI21X1TS \add_x_19_1/U173  ( .A0(\add_x_19_1/n146 ), .A1(\add_x_19_1/n213 ), 
        .B0(\add_x_19_1/n143 ), .Y(\add_x_19_1/n141 ) );
  OAI21X1TS \add_x_19_1/U181  ( .A0(\add_x_19_1/n156 ), .A1(\add_x_19_1/n147 ), 
        .B0(\add_x_19_1/n148 ), .Y(\add_x_19_1/n146 ) );
  OAI21X1TS \add_x_19_1/U156  ( .A0(\add_x_19_1/n133 ), .A1(\add_x_19_1/n131 ), 
        .B0(\add_x_19_1/n132 ), .Y(\add_x_19_1/n130 ) );
  OAI21X1TS \add_x_19_1/U142  ( .A0(\add_x_19_1/n125 ), .A1(\add_x_19_1/n123 ), 
        .B0(\add_x_19_1/n124 ), .Y(\add_x_19_1/n122 ) );
  AOI21X1TS \add_x_19_1/U148  ( .A0(\add_x_19_1/n134 ), .A1(\add_x_19_1/n126 ), 
        .B0(\add_x_19_1/n127 ), .Y(\add_x_19_1/n125 ) );
  OAI21X1TS \add_x_19_1/U163  ( .A0(\add_x_19_1/n156 ), .A1(\add_x_19_1/n135 ), 
        .B0(\add_x_19_1/n136 ), .Y(\add_x_19_1/n134 ) );
  OAI21X1TS \add_x_19_1/U90  ( .A0(\add_x_19_1/n91 ), .A1(\add_x_19_1/n89 ), 
        .B0(\add_x_19_1/n90 ), .Y(\add_x_19_1/n88 ) );
  OAI21X1TS \add_x_19_1/U31  ( .A0(\add_x_19_1/n68 ), .A1(\add_x_19_1/n51 ), 
        .B0(\add_x_19_1/n52 ), .Y(\add_x_19_1/n50 ) );
  OAI21X1TS \add_x_19_1/U55  ( .A0(\add_x_19_1/n68 ), .A1(\add_x_19_1/n66 ), 
        .B0(\add_x_19_1/n67 ), .Y(\add_x_19_1/n65 ) );
  NOR2X1TS \add_x_19_1/U10  ( .A(n1849), .B(n2456), .Y(\add_x_19_1/n36 ) );
  OAI21X1TS \add_x_19_1/U25  ( .A0(\add_x_19_1/n52 ), .A1(\add_x_19_1/n48 ), 
        .B0(\add_x_19_1/n49 ), .Y(\add_x_19_1/n47 ) );
  AOI21X1TS \add_x_19_1/U33  ( .A0(\add_x_19_1/n53 ), .A1(\add_x_19_1/n62 ), 
        .B0(\add_x_19_1/n54 ), .Y(\add_x_19_1/n52 ) );
  OAI21X1TS \add_x_19_1/U35  ( .A0(\add_x_19_1/n55 ), .A1(\add_x_19_1/n59 ), 
        .B0(\add_x_19_1/n56 ), .Y(\add_x_19_1/n54 ) );
  OAI21X1TS \add_x_19_1/U49  ( .A0(\add_x_19_1/n63 ), .A1(\add_x_19_1/n67 ), 
        .B0(\add_x_19_1/n64 ), .Y(\add_x_19_1/n62 ) );
  AOI21X1TS \add_x_19_1/U68  ( .A0(\add_x_19_1/n76 ), .A1(\add_x_19_1/n85 ), 
        .B0(\add_x_19_1/n77 ), .Y(\add_x_19_1/n75 ) );
  OAI21X1TS \add_x_19_1/U84  ( .A0(\add_x_19_1/n86 ), .A1(\add_x_19_1/n90 ), 
        .B0(\add_x_19_1/n87 ), .Y(\add_x_19_1/n85 ) );
  OAI21X1TS \add_x_19_1/U101  ( .A0(\add_x_19_1/n97 ), .A1(\add_x_19_1/n101 ), 
        .B0(\add_x_19_1/n98 ), .Y(\add_x_19_1/n96 ) );
  NOR2X1TS \add_x_19_1/U34  ( .A(\add_x_19_1/n58 ), .B(\add_x_19_1/n55 ), .Y(
        \add_x_19_1/n53 ) );
  NOR2X1TS \add_x_19_1/U48  ( .A(\add_x_19_1/n66 ), .B(\add_x_19_1/n63 ), .Y(
        \add_x_19_1/n61 ) );
  NOR2X1TS \add_x_19_1/U65  ( .A(\add_x_19_1/n93 ), .B(\add_x_19_1/n74 ), .Y(
        \add_x_19_1/n72 ) );
  NOR2X1TS \add_x_19_1/U69  ( .A(\add_x_19_1/n81 ), .B(\add_x_19_1/n78 ), .Y(
        \add_x_19_1/n76 ) );
  NOR2X1TS \add_x_19_1/U83  ( .A(\add_x_19_1/n89 ), .B(\add_x_19_1/n86 ), .Y(
        \add_x_19_1/n84 ) );
  NOR2X1TS \add_x_19_1/U100  ( .A(\add_x_19_1/n100 ), .B(\add_x_19_1/n97 ), 
        .Y(\add_x_19_1/n95 ) );
  OAI21X1TS \add_x_19_1/U150  ( .A0(\add_x_19_1/n128 ), .A1(\add_x_19_1/n132 ), 
        .B0(\add_x_19_1/n129 ), .Y(\add_x_19_1/n127 ) );
  NOR2X1TS \add_x_19_1/U139  ( .A(\addr_calc/fft_write_calc/count[15] ), .B(
        n2475), .Y(\add_x_19_1/n120 ) );
  NOR2X1TS \add_x_19_1/U149  ( .A(\add_x_19_1/n131 ), .B(\add_x_19_1/n128 ), 
        .Y(\add_x_19_1/n126 ) );
  NOR2X1TS \add_x_19_1/U184  ( .A(\add_x_19_1/n154 ), .B(\add_x_19_1/n151 ), 
        .Y(\add_x_19_1/n149 ) );
  NOR2X1TS \add_x_19_1/U249  ( .A(\addr_calc/fft_write_calc/count[1] ), .B(
        n2454), .Y(\add_x_19_1/n188 ) );
  XOR2X1TS \add_x_19_1/U213  ( .A(\add_x_19_1/n172 ), .B(\add_x_19_1/n27 ), 
        .Y(\addr_calc/fft_write_addr[5] ) );
  XOR2X1TS \add_x_19_1/U161  ( .A(\add_x_19_1/n141 ), .B(\add_x_19_1/n21 ), 
        .Y(\addr_calc/fft_write_addr[11] ) );
  NAND2X1TS \add_x_19_1/U11  ( .A(\addr_calc/fft_write_calc/count[30] ), .B(
        n2458), .Y(\add_x_19_1/n37 ) );
  NAND2X1TS \add_x_19_1/U19  ( .A(\addr_calc/fft_write_calc/count[29] ), .B(
        n2388), .Y(\add_x_19_1/n42 ) );
  NAND2X1TS \add_x_19_1/U29  ( .A(n2557), .B(n2386), .Y(\add_x_19_1/n49 ) );
  NAND2X1TS \add_x_19_1/U39  ( .A(n1913), .B(n2500), .Y(\add_x_19_1/n56 ) );
  NAND2X1TS \add_x_19_1/U45  ( .A(\addr_calc/fft_write_calc/count[26] ), .B(
        n2378), .Y(\add_x_19_1/n59 ) );
  NAND2X1TS \add_x_19_1/U53  ( .A(n1915), .B(n2493), .Y(\add_x_19_1/n64 ) );
  NAND2X1TS \add_x_19_1/U74  ( .A(\addr_calc/fft_write_calc/count[23] ), .B(
        n2469), .Y(\add_x_19_1/n79 ) );
  NAND2X1TS \add_x_19_1/U80  ( .A(n2014), .B(n2464), .Y(\add_x_19_1/n82 ) );
  NAND2X1TS \add_x_19_1/U88  ( .A(n1918), .B(n2450), .Y(\add_x_19_1/n87 ) );
  NAND2X1TS \add_x_19_1/U94  ( .A(n2017), .B(n2441), .Y(\add_x_19_1/n90 ) );
  NAND2X1TS \add_x_19_1/U105  ( .A(n1922), .B(n2488), .Y(\add_x_19_1/n98 ) );
  NAND2X1TS \add_x_19_1/U111  ( .A(n2020), .B(n2433), .Y(\add_x_19_1/n101 ) );
  NAND2X1TS \add_x_19_1/U119  ( .A(\addr_calc/fft_write_calc/count[17] ), .B(
        n2479), .Y(\add_x_19_1/n106 ) );
  NOR2X1TS \add_x_19_1/U52  ( .A(n1915), .B(n2493), .Y(\add_x_19_1/n63 ) );
  NOR2X1TS \add_x_19_1/U58  ( .A(n2011), .B(n2460), .Y(\add_x_19_1/n66 ) );
  NOR2X1TS \add_x_19_1/U79  ( .A(n2014), .B(n2464), .Y(\add_x_19_1/n81 ) );
  NOR2X1TS \add_x_19_1/U87  ( .A(n1918), .B(n2448), .Y(\add_x_19_1/n86 ) );
  NOR2X1TS \add_x_19_1/U93  ( .A(n2017), .B(n2440), .Y(\add_x_19_1/n89 ) );
  NOR2X1TS \add_x_19_1/U104  ( .A(n1922), .B(n2487), .Y(\add_x_19_1/n97 ) );
  NOR2X1TS \add_x_19_1/U110  ( .A(n2020), .B(n2432), .Y(\add_x_19_1/n100 ) );
  NOR2X1TS \add_x_19_1/U118  ( .A(\addr_calc/fft_write_calc/count[17] ), .B(
        n2480), .Y(\add_x_19_1/n105 ) );
  NAND2X1TS \add_x_19_1/U140  ( .A(\addr_calc/fft_write_calc/count[15] ), .B(
        n2477), .Y(\add_x_19_1/n121 ) );
  NAND2X1TS \add_x_19_1/U146  ( .A(n2021), .B(n2424), .Y(\add_x_19_1/n124 ) );
  NAND2X1TS \add_x_19_1/U154  ( .A(\addr_calc/fft_write_calc/count[13] ), .B(
        n2417), .Y(\add_x_19_1/n129 ) );
  NAND2X1TS \add_x_19_1/U160  ( .A(\addr_calc/fft_write_calc/count[12] ), .B(
        n2408), .Y(\add_x_19_1/n132 ) );
  NAND2X1TS \add_x_19_1/U179  ( .A(\addr_calc/fft_write_calc/count[10] ), .B(
        n2412), .Y(\add_x_19_1/n145 ) );
  NAND2X1TS \add_x_19_1/U189  ( .A(\addr_calc/fft_write_calc/count[9] ), .B(
        n2496), .Y(\add_x_19_1/n152 ) );
  NOR2X1TS \add_x_19_1/U153  ( .A(\addr_calc/fft_write_calc/count[13] ), .B(
        n2417), .Y(\add_x_19_1/n128 ) );
  NOR2X1TS \add_x_19_1/U159  ( .A(\addr_calc/fft_write_calc/count[12] ), .B(
        n2408), .Y(\add_x_19_1/n131 ) );
  NOR2X1TS \add_x_19_1/U194  ( .A(\addr_calc/fft_write_calc/count[8] ), .B(
        n2472), .Y(\add_x_19_1/n154 ) );
  NAND2X1TS \add_x_19_1/U206  ( .A(\addr_calc/fft_write_calc/count[7] ), .B(
        n2421), .Y(\add_x_19_1/n163 ) );
  NAND2X1TS \add_x_19_1/U212  ( .A(n2030), .B(n2428), .Y(\add_x_19_1/n166 ) );
  NAND2X1TS \add_x_19_1/U228  ( .A(\addr_calc/fft_write_calc/count[4] ), .B(
        n2397), .Y(\add_x_19_1/n176 ) );
  NOR2X1TS \add_x_19_1/U227  ( .A(\addr_calc/fft_write_calc/count[4] ), .B(
        n2397), .Y(\add_x_19_1/n175 ) );
  NAND2X1TS \add_x_19_1/U237  ( .A(\addr_calc/fft_write_calc/count[3] ), .B(
        n2436), .Y(\add_x_19_1/n182 ) );
  NAND2X1TS \add_x_19_1/U243  ( .A(\addr_calc/fft_write_calc/count[2] ), .B(
        n2444), .Y(\add_x_19_1/n185 ) );
  NAND2X1TS \add_x_19_1/U250  ( .A(\addr_calc/fft_write_calc/count[1] ), .B(
        n2452), .Y(\add_x_19_1/n189 ) );
  NOR2X1TS \add_x_19_1/U242  ( .A(\addr_calc/fft_write_calc/count[2] ), .B(
        n2446), .Y(\add_x_19_1/n184 ) );
  XNOR2X1TS \add_x_19_1/U221  ( .A(\add_x_19_1/n177 ), .B(\add_x_19_1/n28 ), 
        .Y(\addr_calc/fft_write_addr[4] ) );
  NAND2X1TS \add_x_19_1/U225  ( .A(\add_x_19_1/n219 ), .B(\add_x_19_1/n176 ), 
        .Y(\add_x_19_1/n28 ) );
  NAND2X1TS \add_x_19_1/U168  ( .A(\add_x_19_1/n212 ), .B(\add_x_19_1/n140 ), 
        .Y(\add_x_19_1/n21 ) );
  XNOR2X1TS \add_x_19_1/U147  ( .A(\add_x_19_1/n130 ), .B(\add_x_19_1/n19 ), 
        .Y(\addr_calc/fft_write_addr[13] ) );
  NAND2X1TS \add_x_19_1/U151  ( .A(\add_x_19_1/n210 ), .B(\add_x_19_1/n129 ), 
        .Y(\add_x_19_1/n19 ) );
  NAND2X1TS \add_x_19_1/U137  ( .A(\add_x_19_1/n208 ), .B(\add_x_19_1/n121 ), 
        .Y(\add_x_19_1/n17 ) );
  XNOR2X1TS \add_x_19_1/U12  ( .A(\add_x_19_1/n3 ), .B(\add_x_19_1/n43 ), .Y(
        \addr_calc/fft_write_addr[29] ) );
  NAND2X1TS \add_x_19_1/U16  ( .A(n2632), .B(\add_x_19_1/n42 ), .Y(
        \add_x_19_1/n3 ) );
  NAND2X1TS \add_x_19_1/U85  ( .A(\add_x_19_1/n202 ), .B(\add_x_19_1/n87 ), 
        .Y(\add_x_19_1/n11 ) );
  NAND2X1TS \add_x_19_1/U26  ( .A(\add_x_19_1/n195 ), .B(\add_x_19_1/n49 ), 
        .Y(\add_x_19_1/n4 ) );
  NAND2X1TS \add_x_19_1/U50  ( .A(\add_x_19_1/n198 ), .B(\add_x_19_1/n64 ), 
        .Y(\add_x_19_1/n7 ) );
  NAND2X1TS \add_x_19_1/U22  ( .A(\add_x_19_1/n72 ), .B(\add_x_19_1/n46 ), .Y(
        \add_x_19_1/n44 ) );
  NAND2X1TS \add_x_19_1/U32  ( .A(\add_x_19_1/n61 ), .B(\add_x_19_1/n53 ), .Y(
        \add_x_19_1/n51 ) );
  NAND2X1TS \add_x_19_1/U67  ( .A(\add_x_19_1/n84 ), .B(\add_x_19_1/n76 ), .Y(
        \add_x_19_1/n74 ) );
  NAND2X1TS \add_x_19_1/U98  ( .A(\add_x_19_1/n103 ), .B(\add_x_19_1/n95 ), 
        .Y(\add_x_19_1/n93 ) );
  NAND2X1TS \add_x_19_1/U171  ( .A(n1667), .B(n2406), .Y(\add_x_19_1/n140 ) );
  NAND2X1TS \add_x_19_1/U133  ( .A(\add_x_19_1/n126 ), .B(\add_x_19_1/n118 ), 
        .Y(\add_x_19_1/n116 ) );
  NAND2X1TS \add_x_19_1/U164  ( .A(\add_x_19_1/n149 ), .B(\add_x_19_1/n137 ), 
        .Y(\add_x_19_1/n135 ) );
  NOR2X2TS \add_x_19_3/U118  ( .A(n1886), .B(n2480), .Y(\add_x_19_3/n105 ) );
  NOR2X1TS \add_x_19_3/U236  ( .A(\addr_calc/fir_write_calc/count[3] ), .B(
        n2438), .Y(\add_x_19_3/n181 ) );
  NOR2X1TS \add_x_19_3/U219  ( .A(\addr_calc/fir_write_calc/count[5] ), .B(
        n2485), .Y(\add_x_19_3/n170 ) );
  OAI21X1TS \add_x_19_3/U70  ( .A0(\add_x_19_3/n78 ), .A1(\add_x_19_3/n82 ), 
        .B0(\add_x_19_3/n79 ), .Y(\add_x_19_3/n77 ) );
  XOR2X1TS \add_x_19_3/U238  ( .A(\add_x_19_3/n186 ), .B(\add_x_19_3/n30 ), 
        .Y(\addr_calc/fir_write_addr[2] ) );
  AOI21X1TS \add_x_19_3/U222  ( .A0(\add_x_19_3/n177 ), .A1(\add_x_19_3/n219 ), 
        .B0(\add_x_19_3/n174 ), .Y(\add_x_19_3/n172 ) );
  AOI21X1TS \add_x_19_3/U214  ( .A0(\add_x_19_3/n177 ), .A1(\add_x_19_3/n168 ), 
        .B0(\add_x_19_3/n169 ), .Y(\add_x_19_3/n167 ) );
  XOR2X1TS \add_x_19_3/U190  ( .A(\add_x_19_3/n156 ), .B(\add_x_19_3/n24 ), 
        .Y(\addr_calc/fir_write_addr[8] ) );
  OAI21X1TS \add_x_19_3/U181  ( .A0(\add_x_19_3/n156 ), .A1(\add_x_19_3/n147 ), 
        .B0(\add_x_19_3/n148 ), .Y(\add_x_19_3/n146 ) );
  OAI21X1TS \add_x_19_3/U142  ( .A0(\add_x_19_3/n125 ), .A1(\add_x_19_3/n123 ), 
        .B0(\add_x_19_3/n124 ), .Y(\add_x_19_3/n122 ) );
  AOI21X1TS \add_x_19_3/U148  ( .A0(\add_x_19_3/n134 ), .A1(\add_x_19_3/n126 ), 
        .B0(\add_x_19_3/n127 ), .Y(\add_x_19_3/n125 ) );
  OAI21X1TS \add_x_19_3/U163  ( .A0(\add_x_19_3/n156 ), .A1(\add_x_19_3/n135 ), 
        .B0(\add_x_19_3/n136 ), .Y(\add_x_19_3/n134 ) );
  OAI21X1TS \add_x_19_3/U107  ( .A0(\add_x_19_3/n102 ), .A1(\add_x_19_3/n100 ), 
        .B0(\add_x_19_3/n101 ), .Y(\add_x_19_3/n99 ) );
  AOI21X1TS \add_x_19_3/U113  ( .A0(n1676), .A1(\add_x_19_3/n103 ), .B0(
        \add_x_19_3/n104 ), .Y(\add_x_19_3/n102 ) );
  OAI21X1TS \add_x_19_3/U90  ( .A0(\add_x_19_3/n91 ), .A1(\add_x_19_3/n89 ), 
        .B0(\add_x_19_3/n90 ), .Y(\add_x_19_3/n88 ) );
  NOR2X1TS \add_x_19_3/U10  ( .A(\addr_calc/fir_write_calc/count[30] ), .B(
        n2456), .Y(\add_x_19_3/n36 ) );
  OAI21X1TS \add_x_19_3/U25  ( .A0(\add_x_19_3/n52 ), .A1(\add_x_19_3/n48 ), 
        .B0(\add_x_19_3/n49 ), .Y(\add_x_19_3/n47 ) );
  OAI21X1TS \add_x_19_3/U35  ( .A0(\add_x_19_3/n55 ), .A1(\add_x_19_3/n59 ), 
        .B0(\add_x_19_3/n56 ), .Y(\add_x_19_3/n54 ) );
  NOR2X1TS \add_x_19_3/U28  ( .A(\addr_calc/fir_write_calc/count[28] ), .B(
        n2386), .Y(\add_x_19_3/n48 ) );
  OAI21X1TS \add_x_19_3/U49  ( .A0(\add_x_19_3/n63 ), .A1(\add_x_19_3/n67 ), 
        .B0(\add_x_19_3/n64 ), .Y(\add_x_19_3/n62 ) );
  NOR2X1TS \add_x_19_3/U48  ( .A(\add_x_19_3/n66 ), .B(\add_x_19_3/n63 ), .Y(
        \add_x_19_3/n61 ) );
  AOI21X1TS \add_x_19_3/U68  ( .A0(\add_x_19_3/n76 ), .A1(\add_x_19_3/n85 ), 
        .B0(\add_x_19_3/n77 ), .Y(\add_x_19_3/n75 ) );
  OAI21X1TS \add_x_19_3/U84  ( .A0(\add_x_19_3/n86 ), .A1(\add_x_19_3/n90 ), 
        .B0(\add_x_19_3/n87 ), .Y(\add_x_19_3/n85 ) );
  OAI21X1TS \add_x_19_3/U101  ( .A0(\add_x_19_3/n97 ), .A1(\add_x_19_3/n101 ), 
        .B0(\add_x_19_3/n98 ), .Y(\add_x_19_3/n96 ) );
  NOR2X1TS \add_x_19_3/U69  ( .A(\add_x_19_3/n81 ), .B(\add_x_19_3/n78 ), .Y(
        \add_x_19_3/n76 ) );
  NOR2X1TS \add_x_19_3/U83  ( .A(\add_x_19_3/n89 ), .B(\add_x_19_3/n86 ), .Y(
        \add_x_19_3/n84 ) );
  NOR2X1TS \add_x_19_3/U100  ( .A(\add_x_19_3/n100 ), .B(\add_x_19_3/n97 ), 
        .Y(\add_x_19_3/n95 ) );
  NOR2X1TS \add_x_19_3/U114  ( .A(\add_x_19_3/n110 ), .B(\add_x_19_3/n105 ), 
        .Y(\add_x_19_3/n103 ) );
  NOR2X1TS \add_x_19_3/U166  ( .A(\add_x_19_3/n144 ), .B(\add_x_19_3/n139 ), 
        .Y(\add_x_19_3/n137 ) );
  NOR2X1TS \add_x_19_3/U170  ( .A(\addr_calc/fir_write_calc/count[11] ), .B(
        n2404), .Y(\add_x_19_3/n139 ) );
  NOR2X1TS \add_x_19_3/U184  ( .A(\add_x_19_3/n154 ), .B(\add_x_19_3/n151 ), 
        .Y(\add_x_19_3/n149 ) );
  NOR2X1TS \add_x_19_3/U215  ( .A(\add_x_19_3/n175 ), .B(\add_x_19_3/n170 ), 
        .Y(\add_x_19_3/n168 ) );
  NOR2X1TS \add_x_19_3/U249  ( .A(\addr_calc/fir_write_calc/count[1] ), .B(
        n2454), .Y(\add_x_19_3/n188 ) );
  XOR2X1TS \add_x_19_3/U213  ( .A(\add_x_19_3/n172 ), .B(\add_x_19_3/n27 ), 
        .Y(\addr_calc/fir_write_addr[5] ) );
  XOR2X1TS \add_x_19_3/U207  ( .A(\add_x_19_3/n167 ), .B(\add_x_19_3/n26 ), 
        .Y(\addr_calc/fir_write_addr[6] ) );
  XOR2X1TS \add_x_19_3/U141  ( .A(\add_x_19_3/n125 ), .B(\add_x_19_3/n18 ), 
        .Y(\addr_calc/fir_write_addr[14] ) );
  NAND2X1TS \add_x_19_3/U11  ( .A(n1836), .B(n2458), .Y(\add_x_19_3/n37 ) );
  NAND2X1TS \add_x_19_3/U19  ( .A(\addr_calc/fir_write_calc/count[29] ), .B(
        n2390), .Y(\add_x_19_3/n42 ) );
  NAND2X1TS \add_x_19_3/U29  ( .A(n1896), .B(n2386), .Y(\add_x_19_3/n49 ) );
  NAND2X1TS \add_x_19_3/U39  ( .A(n1835), .B(n2499), .Y(\add_x_19_3/n56 ) );
  NAND2X1TS \add_x_19_3/U45  ( .A(\addr_calc/fir_write_calc/count[26] ), .B(
        n2377), .Y(\add_x_19_3/n59 ) );
  NAND2X1TS \add_x_19_3/U53  ( .A(\addr_calc/fir_write_calc/count[25] ), .B(
        n2492), .Y(\add_x_19_3/n64 ) );
  NAND2X1TS \add_x_19_3/U59  ( .A(\addr_calc/fir_write_calc/count[24] ), .B(
        n2461), .Y(\add_x_19_3/n67 ) );
  NAND2X1TS \add_x_19_3/U74  ( .A(\addr_calc/fir_write_calc/count[23] ), .B(
        n2469), .Y(\add_x_19_3/n79 ) );
  NAND2X1TS \add_x_19_3/U80  ( .A(\addr_calc/fir_write_calc/count[22] ), .B(
        n2466), .Y(\add_x_19_3/n82 ) );
  NAND2X1TS \add_x_19_3/U88  ( .A(n1892), .B(n2450), .Y(\add_x_19_3/n87 ) );
  NAND2X1TS \add_x_19_3/U94  ( .A(n2009), .B(n2442), .Y(\add_x_19_3/n90 ) );
  NAND2X1TS \add_x_19_3/U105  ( .A(n1670), .B(n2488), .Y(\add_x_19_3/n98 ) );
  NAND2X1TS \add_x_19_3/U111  ( .A(\addr_calc/fir_write_calc/count[18] ), .B(
        n2434), .Y(\add_x_19_3/n101 ) );
  NOR2X1TS \add_x_19_3/U79  ( .A(n1668), .B(n2465), .Y(\add_x_19_3/n81 ) );
  NOR2X1TS \add_x_19_3/U93  ( .A(n1669), .B(n2442), .Y(\add_x_19_3/n89 ) );
  NOR2X1TS \add_x_19_3/U110  ( .A(n2006), .B(n2434), .Y(\add_x_19_3/n100 ) );
  NAND2X1TS \add_x_19_3/U140  ( .A(n1883), .B(n2476), .Y(\add_x_19_3/n121 ) );
  NAND2X1TS \add_x_19_3/U146  ( .A(n2003), .B(n2425), .Y(\add_x_19_3/n124 ) );
  NAND2X1TS \add_x_19_3/U154  ( .A(\addr_calc/fir_write_calc/count[13] ), .B(
        n2418), .Y(\add_x_19_3/n129 ) );
  NAND2X1TS \add_x_19_3/U179  ( .A(\addr_calc/fir_write_calc/count[10] ), .B(
        n2414), .Y(\add_x_19_3/n145 ) );
  NAND2X1TS \add_x_19_3/U189  ( .A(\addr_calc/fir_write_calc/count[9] ), .B(
        n2496), .Y(\add_x_19_3/n152 ) );
  NOR2X1TS \add_x_19_3/U153  ( .A(\addr_calc/fir_write_calc/count[13] ), .B(
        n2418), .Y(\add_x_19_3/n128 ) );
  NOR2X1TS \add_x_19_3/U178  ( .A(\addr_calc/fir_write_calc/count[10] ), .B(
        n2413), .Y(\add_x_19_3/n144 ) );
  NOR2X1TS \add_x_19_3/U188  ( .A(\addr_calc/fir_write_calc/count[9] ), .B(
        n2495), .Y(\add_x_19_3/n151 ) );
  NOR2X1TS \add_x_19_3/U194  ( .A(n1995), .B(n2473), .Y(\add_x_19_3/n154 ) );
  NAND2X1TS \add_x_19_3/U206  ( .A(\addr_calc/fir_write_calc/count[7] ), .B(
        n2420), .Y(\add_x_19_3/n163 ) );
  NAND2X1TS \add_x_19_3/U212  ( .A(n1992), .B(n2430), .Y(\add_x_19_3/n166 ) );
  NAND2X1TS \add_x_19_3/U228  ( .A(n1865), .B(n2396), .Y(\add_x_19_3/n176 ) );
  NOR2X1TS \add_x_19_3/U227  ( .A(n1865), .B(n2397), .Y(\add_x_19_3/n175 ) );
  NAND2X1TS \add_x_19_3/U237  ( .A(\addr_calc/fir_write_calc/count[3] ), .B(
        n2437), .Y(\add_x_19_3/n182 ) );
  NAND2X1TS \add_x_19_3/U250  ( .A(n2452), .B(
        \addr_calc/fir_write_calc/count[1] ), .Y(\add_x_19_3/n189 ) );
  NAND2X1TS \add_x_19_3/U240  ( .A(\add_x_19_3/n221 ), .B(\add_x_19_3/n185 ), 
        .Y(\add_x_19_3/n30 ) );
  XNOR2X1TS \add_x_19_3/U221  ( .A(\add_x_19_3/n177 ), .B(\add_x_19_3/n28 ), 
        .Y(\addr_calc/fir_write_addr[4] ) );
  NAND2X1TS \add_x_19_3/U225  ( .A(\add_x_19_3/n219 ), .B(\add_x_19_3/n176 ), 
        .Y(\add_x_19_3/n28 ) );
  NAND2X1TS \add_x_19_3/U217  ( .A(\add_x_19_3/n218 ), .B(\add_x_19_3/n171 ), 
        .Y(\add_x_19_3/n27 ) );
  NAND2X1TS \add_x_19_3/U209  ( .A(\add_x_19_3/n217 ), .B(\add_x_19_3/n166 ), 
        .Y(\add_x_19_3/n26 ) );
  NAND2X1TS \add_x_19_3/U192  ( .A(\add_x_19_3/n215 ), .B(\add_x_19_3/n155 ), 
        .Y(\add_x_19_3/n24 ) );
  XNOR2X1TS \add_x_19_3/U172  ( .A(\add_x_19_3/n146 ), .B(\add_x_19_3/n22 ), 
        .Y(\addr_calc/fir_write_addr[10] ) );
  NAND2X1TS \add_x_19_3/U176  ( .A(\add_x_19_3/n213 ), .B(\add_x_19_3/n145 ), 
        .Y(\add_x_19_3/n22 ) );
  NAND2X1TS \add_x_19_3/U143  ( .A(n1545), .B(\add_x_19_3/n124 ), .Y(
        \add_x_19_3/n18 ) );
  XNOR2X1TS \add_x_19_3/U128  ( .A(\add_x_19_3/n122 ), .B(\add_x_19_3/n17 ), 
        .Y(\addr_calc/fir_write_addr[15] ) );
  NAND2X1TS \add_x_19_3/U137  ( .A(\add_x_19_3/n208 ), .B(\add_x_19_3/n121 ), 
        .Y(\add_x_19_3/n17 ) );
  XNOR2X1TS \add_x_19_3/U95  ( .A(\add_x_19_3/n99 ), .B(\add_x_19_3/n13 ), .Y(
        \addr_calc/fir_write_addr[19] ) );
  NAND2X1TS \add_x_19_3/U102  ( .A(\add_x_19_3/n204 ), .B(\add_x_19_3/n98 ), 
        .Y(\add_x_19_3/n13 ) );
  XNOR2X1TS \add_x_19_3/U81  ( .A(\add_x_19_3/n88 ), .B(\add_x_19_3/n11 ), .Y(
        \addr_calc/fir_write_addr[21] ) );
  NAND2X1TS \add_x_19_3/U85  ( .A(\add_x_19_3/n202 ), .B(\add_x_19_3/n87 ), 
        .Y(\add_x_19_3/n11 ) );
  NAND2X1TS \add_x_19_3/U26  ( .A(\add_x_19_3/n195 ), .B(\add_x_19_3/n49 ), 
        .Y(\add_x_19_3/n4 ) );
  XNOR2X1TS \add_x_19_3/U46  ( .A(\add_x_19_3/n65 ), .B(\add_x_19_3/n7 ), .Y(
        \addr_calc/fir_write_addr[25] ) );
  NAND2X1TS \add_x_19_3/U50  ( .A(\add_x_19_3/n198 ), .B(\add_x_19_3/n64 ), 
        .Y(\add_x_19_3/n7 ) );
  NAND2X1TS \add_x_19_3/U119  ( .A(n1886), .B(n2481), .Y(\add_x_19_3/n106 ) );
  NAND2X1TS \add_x_19_3/U67  ( .A(\add_x_19_3/n84 ), .B(\add_x_19_3/n76 ), .Y(
        \add_x_19_3/n74 ) );
  NAND2X1TS \add_x_19_3/U98  ( .A(\add_x_19_3/n103 ), .B(\add_x_19_3/n95 ), 
        .Y(\add_x_19_3/n93 ) );
  NAND2X1TS \add_x_19_3/U171  ( .A(\addr_calc/fir_write_calc/count[11] ), .B(
        n2405), .Y(\add_x_19_3/n140 ) );
  NAND2X1TS \add_x_19_3/U164  ( .A(\add_x_19_3/n149 ), .B(\add_x_19_3/n137 ), 
        .Y(\add_x_19_3/n135 ) );
  NAND2X1TS \add_x_19_3/U220  ( .A(\addr_calc/fir_write_calc/count[5] ), .B(
        n2483), .Y(\add_x_19_3/n171 ) );
  NOR2X1TS \add_x_19_5/U236  ( .A(n1933), .B(n2437), .Y(\add_x_19_5/n181 ) );
  OAI21X2TS \add_x_19_5/U198  ( .A0(\add_x_19_5/n178 ), .A1(\add_x_19_5/n158 ), 
        .B0(\add_x_19_5/n159 ), .Y(\add_x_19_5/n157 ) );
  NAND2X1TS \add_x_19_5/U255  ( .A(\addr_calc/iir_write_calc/count[0] ), .B(
        n2392), .Y(\add_x_19_5/n191 ) );
  XOR2X1TS \add_x_19_5/U244  ( .A(\add_x_19_5/n31 ), .B(\add_x_19_5/n191 ), 
        .Y(\addr_calc/iir_write_addr[1] ) );
  AOI21X1TS \add_x_19_5/U214  ( .A0(n1818), .A1(\add_x_19_5/n168 ), .B0(
        \add_x_19_5/n169 ), .Y(\add_x_19_5/n167 ) );
  OAI21X1TS \add_x_19_5/U191  ( .A0(\add_x_19_5/n156 ), .A1(\add_x_19_5/n154 ), 
        .B0(\add_x_19_5/n155 ), .Y(\add_x_19_5/n153 ) );
  OAI21X1TS \add_x_19_5/U181  ( .A0(\add_x_19_5/n156 ), .A1(\add_x_19_5/n147 ), 
        .B0(\add_x_19_5/n148 ), .Y(\add_x_19_5/n146 ) );
  OAI21X1TS \add_x_19_5/U156  ( .A0(\add_x_19_5/n133 ), .A1(\add_x_19_5/n131 ), 
        .B0(\add_x_19_5/n132 ), .Y(\add_x_19_5/n130 ) );
  AOI21X1TS \add_x_19_5/U121  ( .A0(\add_x_19_5/n112 ), .A1(\add_x_19_5/n207 ), 
        .B0(\add_x_19_5/n109 ), .Y(\add_x_19_5/n107 ) );
  OAI21X1TS \add_x_19_5/U90  ( .A0(\add_x_19_5/n91 ), .A1(\add_x_19_5/n89 ), 
        .B0(\add_x_19_5/n90 ), .Y(\add_x_19_5/n88 ) );
  OAI21X1TS \add_x_19_5/U31  ( .A0(\add_x_19_5/n68 ), .A1(\add_x_19_5/n51 ), 
        .B0(\add_x_19_5/n52 ), .Y(\add_x_19_5/n50 ) );
  OAI21X1TS \add_x_19_5/U55  ( .A0(\add_x_19_5/n68 ), .A1(\add_x_19_5/n66 ), 
        .B0(\add_x_19_5/n67 ), .Y(\add_x_19_5/n65 ) );
  NOR2X1TS \add_x_19_5/U10  ( .A(\addr_calc/iir_write_calc/count[30] ), .B(
        n2457), .Y(\add_x_19_5/n36 ) );
  OAI21X1TS \add_x_19_5/U49  ( .A0(\add_x_19_5/n63 ), .A1(\add_x_19_5/n67 ), 
        .B0(\add_x_19_5/n64 ), .Y(\add_x_19_5/n62 ) );
  AOI21X1TS \add_x_19_5/U99  ( .A0(\add_x_19_5/n95 ), .A1(\add_x_19_5/n104 ), 
        .B0(\add_x_19_5/n96 ), .Y(\add_x_19_5/n94 ) );
  OAI21X1TS \add_x_19_5/U101  ( .A0(\add_x_19_5/n97 ), .A1(\add_x_19_5/n101 ), 
        .B0(\add_x_19_5/n98 ), .Y(\add_x_19_5/n96 ) );
  NOR2X1TS \add_x_19_5/U28  ( .A(n1974), .B(n2385), .Y(\add_x_19_5/n48 ) );
  NOR2X1TS \add_x_19_5/U34  ( .A(\add_x_19_5/n58 ), .B(\add_x_19_5/n55 ), .Y(
        \add_x_19_5/n53 ) );
  NOR2X1TS \add_x_19_5/U48  ( .A(\add_x_19_5/n66 ), .B(\add_x_19_5/n63 ), .Y(
        \add_x_19_5/n61 ) );
  NOR2X1TS \add_x_19_5/U65  ( .A(\add_x_19_5/n93 ), .B(\add_x_19_5/n74 ), .Y(
        \add_x_19_5/n72 ) );
  NOR2X1TS \add_x_19_5/U83  ( .A(\add_x_19_5/n89 ), .B(\add_x_19_5/n86 ), .Y(
        \add_x_19_5/n84 ) );
  NOR2X1TS \add_x_19_5/U100  ( .A(\add_x_19_5/n100 ), .B(\add_x_19_5/n97 ), 
        .Y(\add_x_19_5/n95 ) );
  OAI21X1TS \add_x_19_5/U150  ( .A0(\add_x_19_5/n128 ), .A1(\add_x_19_5/n132 ), 
        .B0(\add_x_19_5/n129 ), .Y(\add_x_19_5/n127 ) );
  OAI21X1TS \add_x_19_5/U167  ( .A0(\add_x_19_5/n139 ), .A1(\add_x_19_5/n145 ), 
        .B0(\add_x_19_5/n140 ), .Y(\add_x_19_5/n138 ) );
  OAI21X1TS \add_x_19_5/U185  ( .A0(\add_x_19_5/n151 ), .A1(\add_x_19_5/n155 ), 
        .B0(\add_x_19_5/n152 ), .Y(\add_x_19_5/n150 ) );
  NOR2X1TS \add_x_19_5/U139  ( .A(\addr_calc/iir_write_calc/count[15] ), .B(
        n2477), .Y(\add_x_19_5/n120 ) );
  NOR2X1TS \add_x_19_5/U149  ( .A(\add_x_19_5/n131 ), .B(\add_x_19_5/n128 ), 
        .Y(\add_x_19_5/n126 ) );
  NOR2X1TS \add_x_19_5/U166  ( .A(\add_x_19_5/n144 ), .B(\add_x_19_5/n139 ), 
        .Y(\add_x_19_5/n137 ) );
  NOR2X1TS \add_x_19_5/U170  ( .A(\addr_calc/iir_write_calc/count[11] ), .B(
        n2405), .Y(\add_x_19_5/n139 ) );
  NOR2X1TS \add_x_19_5/U184  ( .A(\add_x_19_5/n154 ), .B(\add_x_19_5/n151 ), 
        .Y(\add_x_19_5/n149 ) );
  AOI21X1TS \add_x_19_5/U200  ( .A0(\add_x_19_5/n160 ), .A1(\add_x_19_5/n169 ), 
        .B0(\add_x_19_5/n161 ), .Y(\add_x_19_5/n159 ) );
  OAI21X1TS \add_x_19_5/U202  ( .A0(\add_x_19_5/n162 ), .A1(\add_x_19_5/n166 ), 
        .B0(\add_x_19_5/n163 ), .Y(\add_x_19_5/n161 ) );
  OAI21X1TS \add_x_19_5/U216  ( .A0(\add_x_19_5/n170 ), .A1(\add_x_19_5/n176 ), 
        .B0(\add_x_19_5/n171 ), .Y(\add_x_19_5/n169 ) );
  NOR2X1TS \add_x_19_5/U201  ( .A(\add_x_19_5/n165 ), .B(\add_x_19_5/n162 ), 
        .Y(\add_x_19_5/n160 ) );
  NOR2X1TS \add_x_19_5/U215  ( .A(\add_x_19_5/n175 ), .B(\add_x_19_5/n170 ), 
        .Y(\add_x_19_5/n168 ) );
  AOI21X1TS \add_x_19_5/U231  ( .A0(\add_x_19_5/n179 ), .A1(\add_x_19_5/n187 ), 
        .B0(\add_x_19_5/n180 ), .Y(\add_x_19_5/n178 ) );
  OAI21X1TS \add_x_19_5/U233  ( .A0(\add_x_19_5/n181 ), .A1(\add_x_19_5/n185 ), 
        .B0(\add_x_19_5/n182 ), .Y(\add_x_19_5/n180 ) );
  OAI21X1TS \add_x_19_5/U246  ( .A0(\add_x_19_5/n188 ), .A1(\add_x_19_5/n191 ), 
        .B0(\add_x_19_5/n189 ), .Y(\add_x_19_5/n187 ) );
  NOR2X1TS \add_x_19_5/U249  ( .A(\addr_calc/iir_write_calc/count[1] ), .B(
        n2452), .Y(\add_x_19_5/n188 ) );
  NOR2X1TS \add_x_19_5/U232  ( .A(\add_x_19_5/n184 ), .B(\add_x_19_5/n181 ), 
        .Y(\add_x_19_5/n179 ) );
  XOR2X1TS \add_x_19_5/U112  ( .A(\add_x_19_5/n107 ), .B(\add_x_19_5/n15 ), 
        .Y(\addr_calc/iir_write_addr[17] ) );
  NAND2X1TS \add_x_19_5/U11  ( .A(n1854), .B(n2456), .Y(\add_x_19_5/n37 ) );
  NAND2X1TS \add_x_19_5/U19  ( .A(n1851), .B(n2388), .Y(\add_x_19_5/n42 ) );
  NAND2X1TS \add_x_19_5/U29  ( .A(\addr_calc/iir_write_calc/count[28] ), .B(
        n2384), .Y(\add_x_19_5/n49 ) );
  NAND2X1TS \add_x_19_5/U39  ( .A(\addr_calc/iir_write_calc/count[27] ), .B(
        n2499), .Y(\add_x_19_5/n56 ) );
  NAND2X1TS \add_x_19_5/U45  ( .A(\addr_calc/iir_write_calc/count[26] ), .B(
        n2378), .Y(\add_x_19_5/n59 ) );
  NAND2X1TS \add_x_19_5/U53  ( .A(n1969), .B(n2491), .Y(\add_x_19_5/n64 ) );
  NAND2X1TS \add_x_19_5/U59  ( .A(n2051), .B(n2461), .Y(\add_x_19_5/n67 ) );
  NAND2X1TS \add_x_19_5/U74  ( .A(n1965), .B(n2470), .Y(\add_x_19_5/n79 ) );
  NAND2X1TS \add_x_19_5/U80  ( .A(\addr_calc/iir_write_calc/count[22] ), .B(
        n2465), .Y(\add_x_19_5/n82 ) );
  NAND2X1TS \add_x_19_5/U88  ( .A(n1962), .B(n2449), .Y(\add_x_19_5/n87 ) );
  NAND2X1TS \add_x_19_5/U105  ( .A(n1958), .B(n2489), .Y(\add_x_19_5/n98 ) );
  NAND2X1TS \add_x_19_5/U111  ( .A(\addr_calc/iir_write_calc/count[18] ), .B(
        n2433), .Y(\add_x_19_5/n101 ) );
  NOR2X1TS \add_x_19_5/U52  ( .A(n1969), .B(n2492), .Y(\add_x_19_5/n63 ) );
  NOR2X1TS \add_x_19_5/U58  ( .A(n2051), .B(n2462), .Y(\add_x_19_5/n66 ) );
  NOR2X1TS \add_x_19_5/U87  ( .A(n1962), .B(n2449), .Y(\add_x_19_5/n86 ) );
  NOR2X1TS \add_x_19_5/U93  ( .A(n2048), .B(n2441), .Y(\add_x_19_5/n89 ) );
  NOR2X1TS \add_x_19_5/U110  ( .A(\addr_calc/iir_write_calc/count[18] ), .B(
        n2433), .Y(\add_x_19_5/n100 ) );
  NOR2X1TS \add_x_19_5/U118  ( .A(\addr_calc/iir_write_calc/count[17] ), .B(
        n2480), .Y(\add_x_19_5/n105 ) );
  NOR2X1TS \add_x_19_5/U126  ( .A(\addr_calc/iir_write_calc/count[16] ), .B(
        n2400), .Y(\add_x_19_5/n110 ) );
  NAND2X1TS \add_x_19_5/U140  ( .A(\addr_calc/iir_write_calc/count[15] ), .B(
        n2476), .Y(\add_x_19_5/n121 ) );
  NAND2X1TS \add_x_19_5/U146  ( .A(\addr_calc/iir_write_calc/count[14] ), .B(
        n2426), .Y(\add_x_19_5/n124 ) );
  NAND2X1TS \add_x_19_5/U154  ( .A(\addr_calc/iir_write_calc/count[13] ), .B(
        n2418), .Y(\add_x_19_5/n129 ) );
  NAND2X1TS \add_x_19_5/U160  ( .A(\addr_calc/iir_write_calc/count[12] ), .B(
        n2409), .Y(\add_x_19_5/n132 ) );
  NAND2X1TS \add_x_19_5/U179  ( .A(\addr_calc/iir_write_calc/count[10] ), .B(
        n2414), .Y(\add_x_19_5/n145 ) );
  NAND2X1TS \add_x_19_5/U189  ( .A(\addr_calc/iir_write_calc/count[9] ), .B(
        n1980), .Y(\add_x_19_5/n152 ) );
  NAND2X1TS \add_x_19_5/U195  ( .A(\addr_calc/iir_write_calc/count[8] ), .B(
        n1864), .Y(\add_x_19_5/n155 ) );
  NOR2X1TS \add_x_19_5/U145  ( .A(\addr_calc/iir_write_calc/count[14] ), .B(
        n2425), .Y(\add_x_19_5/n123 ) );
  NOR2X1TS \add_x_19_5/U153  ( .A(\addr_calc/iir_write_calc/count[13] ), .B(
        n2417), .Y(\add_x_19_5/n128 ) );
  NOR2X1TS \add_x_19_5/U159  ( .A(\addr_calc/iir_write_calc/count[12] ), .B(
        n2410), .Y(\add_x_19_5/n131 ) );
  NOR2X1TS \add_x_19_5/U178  ( .A(\addr_calc/iir_write_calc/count[10] ), .B(
        n2414), .Y(\add_x_19_5/n144 ) );
  NOR2X1TS \add_x_19_5/U188  ( .A(\addr_calc/iir_write_calc/count[9] ), .B(
        n2495), .Y(\add_x_19_5/n151 ) );
  NOR2X1TS \add_x_19_5/U194  ( .A(\addr_calc/iir_write_calc/count[8] ), .B(
        n1864), .Y(\add_x_19_5/n154 ) );
  NAND2X1TS \add_x_19_5/U206  ( .A(n1683), .B(n2422), .Y(\add_x_19_5/n163 ) );
  NAND2X1TS \add_x_19_5/U212  ( .A(\addr_calc/iir_write_calc/count[6] ), .B(
        n2429), .Y(\add_x_19_5/n166 ) );
  NAND2X1TS \add_x_19_5/U228  ( .A(\addr_calc/iir_write_calc/count[4] ), .B(
        n2396), .Y(\add_x_19_5/n176 ) );
  NOR2X1TS \add_x_19_5/U211  ( .A(\addr_calc/iir_write_calc/count[6] ), .B(
        n2429), .Y(\add_x_19_5/n165 ) );
  NOR2X1TS \add_x_19_5/U227  ( .A(\addr_calc/iir_write_calc/count[4] ), .B(
        n2398), .Y(\add_x_19_5/n175 ) );
  NAND2X1TS \add_x_19_5/U237  ( .A(n1933), .B(n2437), .Y(\add_x_19_5/n182 ) );
  NAND2X1TS \add_x_19_5/U243  ( .A(\addr_calc/iir_write_calc/count[2] ), .B(
        n2444), .Y(\add_x_19_5/n185 ) );
  NAND2X1TS \add_x_19_5/U250  ( .A(\addr_calc/iir_write_calc/count[1] ), .B(
        n2453), .Y(\add_x_19_5/n189 ) );
  NOR2X1TS \add_x_19_5/U242  ( .A(\addr_calc/iir_write_calc/count[2] ), .B(
        n2445), .Y(\add_x_19_5/n184 ) );
  NAND2X1TS \add_x_19_5/U247  ( .A(\add_x_19_5/n222 ), .B(\add_x_19_5/n189 ), 
        .Y(\add_x_19_5/n31 ) );
  XNOR2X1TS \add_x_19_5/U229  ( .A(\add_x_19_5/n183 ), .B(\add_x_19_5/n29 ), 
        .Y(\addr_calc/iir_write_addr[3] ) );
  NAND2X1TS \add_x_19_5/U234  ( .A(\add_x_19_5/n220 ), .B(\add_x_19_5/n182 ), 
        .Y(\add_x_19_5/n29 ) );
  XNOR2X1TS \add_x_19_5/U221  ( .A(n1818), .B(\add_x_19_5/n28 ), .Y(
        \addr_calc/iir_write_addr[4] ) );
  NAND2X1TS \add_x_19_5/U225  ( .A(\add_x_19_5/n219 ), .B(\add_x_19_5/n176 ), 
        .Y(\add_x_19_5/n28 ) );
  XNOR2X1TS \add_x_19_5/U180  ( .A(\add_x_19_5/n153 ), .B(\add_x_19_5/n23 ), 
        .Y(\addr_calc/iir_write_addr[9] ) );
  NAND2X1TS \add_x_19_5/U186  ( .A(\add_x_19_5/n214 ), .B(\add_x_19_5/n152 ), 
        .Y(\add_x_19_5/n23 ) );
  XNOR2X1TS \add_x_19_5/U172  ( .A(\add_x_19_5/n146 ), .B(\add_x_19_5/n22 ), 
        .Y(\addr_calc/iir_write_addr[10] ) );
  NAND2X1TS \add_x_19_5/U176  ( .A(\add_x_19_5/n213 ), .B(\add_x_19_5/n145 ), 
        .Y(\add_x_19_5/n22 ) );
  XNOR2X1TS \add_x_19_5/U120  ( .A(\add_x_19_5/n112 ), .B(\add_x_19_5/n16 ), 
        .Y(\addr_calc/iir_write_addr[16] ) );
  NAND2X1TS \add_x_19_5/U124  ( .A(\add_x_19_5/n207 ), .B(\add_x_19_5/n111 ), 
        .Y(\add_x_19_5/n16 ) );
  XNOR2X1TS \add_x_19_5/U147  ( .A(\add_x_19_5/n130 ), .B(\add_x_19_5/n19 ), 
        .Y(\addr_calc/iir_write_addr[13] ) );
  NAND2X1TS \add_x_19_5/U151  ( .A(\add_x_19_5/n210 ), .B(\add_x_19_5/n129 ), 
        .Y(\add_x_19_5/n19 ) );
  NAND2X1TS \add_x_19_5/U116  ( .A(\add_x_19_5/n206 ), .B(\add_x_19_5/n106 ), 
        .Y(\add_x_19_5/n15 ) );
  XNOR2X1TS \add_x_19_5/U81  ( .A(\add_x_19_5/n88 ), .B(\add_x_19_5/n11 ), .Y(
        \addr_calc/iir_write_addr[21] ) );
  NAND2X1TS \add_x_19_5/U85  ( .A(\add_x_19_5/n202 ), .B(\add_x_19_5/n87 ), 
        .Y(\add_x_19_5/n11 ) );
  NAND2X1TS \add_x_19_5/U26  ( .A(\add_x_19_5/n195 ), .B(\add_x_19_5/n49 ), 
        .Y(\add_x_19_5/n4 ) );
  NAND2X1TS \add_x_19_5/U50  ( .A(\add_x_19_5/n198 ), .B(\add_x_19_5/n64 ), 
        .Y(\add_x_19_5/n7 ) );
  NAND2X1TS \add_x_19_5/U119  ( .A(\addr_calc/iir_write_calc/count[17] ), .B(
        n2479), .Y(\add_x_19_5/n106 ) );
  NAND2X1TS \add_x_19_5/U32  ( .A(\add_x_19_5/n61 ), .B(\add_x_19_5/n53 ), .Y(
        \add_x_19_5/n51 ) );
  NAND2X1TS \add_x_19_5/U98  ( .A(\add_x_19_5/n103 ), .B(\add_x_19_5/n95 ), 
        .Y(\add_x_19_5/n93 ) );
  NAND2X1TS \add_x_19_5/U171  ( .A(\addr_calc/iir_write_calc/count[11] ), .B(
        n2405), .Y(\add_x_19_5/n140 ) );
  NAND2X1TS \add_x_19_5/U164  ( .A(\add_x_19_5/n149 ), .B(\add_x_19_5/n137 ), 
        .Y(\add_x_19_5/n135 ) );
  NAND2X1TS \add_x_19_5/U220  ( .A(n1686), .B(n2485), .Y(\add_x_19_5/n171 ) );
  NAND2X1TS \add_x_19_5/U199  ( .A(\add_x_19_5/n168 ), .B(\add_x_19_5/n160 ), 
        .Y(\add_x_19_5/n158 ) );
  NOR2X1TS \add_x_19_0/U236  ( .A(\addr_calc/fft_read_calc/count[3] ), .B(
        n2438), .Y(\add_x_19_0/n181 ) );
  NOR2X1TS \add_x_19_0/U219  ( .A(\addr_calc/fft_read_calc/count[5] ), .B(
        n2484), .Y(\add_x_19_0/n170 ) );
  NAND2X1TS \add_x_19_0/U127  ( .A(\addr_calc/fft_read_calc/count[16] ), .B(
        n2402), .Y(\add_x_19_0/n111 ) );
  AOI21X1TS \add_x_19_0/U214  ( .A0(\add_x_19_0/n177 ), .A1(\add_x_19_0/n168 ), 
        .B0(\add_x_19_0/n169 ), .Y(\add_x_19_0/n167 ) );
  XOR2X1TS \add_x_19_0/U190  ( .A(\add_x_19_0/n156 ), .B(\add_x_19_0/n24 ), 
        .Y(\addr_calc/fft_read_addr[8] ) );
  OAI21X1TS \add_x_19_0/U156  ( .A0(\add_x_19_0/n133 ), .A1(\add_x_19_0/n131 ), 
        .B0(\add_x_19_0/n132 ), .Y(\add_x_19_0/n130 ) );
  OAI21X1TS \add_x_19_0/U181  ( .A0(\add_x_19_0/n156 ), .A1(\add_x_19_0/n147 ), 
        .B0(\add_x_19_0/n148 ), .Y(\add_x_19_0/n146 ) );
  OAI21X1TS \add_x_19_0/U142  ( .A0(\add_x_19_0/n125 ), .A1(\add_x_19_0/n123 ), 
        .B0(\add_x_19_0/n124 ), .Y(\add_x_19_0/n122 ) );
  AOI21X1TS \add_x_19_0/U148  ( .A0(\add_x_19_0/n134 ), .A1(\add_x_19_0/n126 ), 
        .B0(\add_x_19_0/n127 ), .Y(\add_x_19_0/n125 ) );
  OAI21X1TS \add_x_19_0/U163  ( .A0(\add_x_19_0/n156 ), .A1(\add_x_19_0/n135 ), 
        .B0(\add_x_19_0/n136 ), .Y(\add_x_19_0/n134 ) );
  AOI21X1TS \add_x_19_0/U121  ( .A0(\add_x_19_0/n112 ), .A1(\add_x_19_0/n207 ), 
        .B0(\add_x_19_0/n109 ), .Y(\add_x_19_0/n107 ) );
  OAI21X1TS \add_x_19_0/U107  ( .A0(\add_x_19_0/n102 ), .A1(\add_x_19_0/n100 ), 
        .B0(\add_x_19_0/n101 ), .Y(\add_x_19_0/n99 ) );
  AOI21X1TS \add_x_19_0/U113  ( .A0(\add_x_19_0/n112 ), .A1(\add_x_19_0/n103 ), 
        .B0(\add_x_19_0/n104 ), .Y(\add_x_19_0/n102 ) );
  OAI21X1TS \add_x_19_0/U90  ( .A0(\add_x_19_0/n91 ), .A1(\add_x_19_0/n89 ), 
        .B0(\add_x_19_0/n90 ), .Y(\add_x_19_0/n88 ) );
  OAI21X1TS \add_x_19_0/U31  ( .A0(\add_x_19_0/n68 ), .A1(\add_x_19_0/n51 ), 
        .B0(\add_x_19_0/n52 ), .Y(\add_x_19_0/n50 ) );
  OAI21X1TS \add_x_19_0/U55  ( .A0(\add_x_19_0/n68 ), .A1(\add_x_19_0/n66 ), 
        .B0(\add_x_19_0/n67 ), .Y(\add_x_19_0/n65 ) );
  NOR2X1TS \add_x_19_0/U10  ( .A(n1859), .B(n2457), .Y(\add_x_19_0/n36 ) );
  AOI21X1TS \add_x_19_0/U23  ( .A0(\add_x_19_0/n73 ), .A1(\add_x_19_0/n46 ), 
        .B0(\add_x_19_0/n47 ), .Y(\add_x_19_0/n45 ) );
  OAI21X1TS \add_x_19_0/U25  ( .A0(\add_x_19_0/n52 ), .A1(\add_x_19_0/n48 ), 
        .B0(\add_x_19_0/n49 ), .Y(\add_x_19_0/n47 ) );
  OAI21X1TS \add_x_19_0/U35  ( .A0(\add_x_19_0/n55 ), .A1(\add_x_19_0/n59 ), 
        .B0(\add_x_19_0/n56 ), .Y(\add_x_19_0/n54 ) );
  OAI21X1TS \add_x_19_0/U49  ( .A0(\add_x_19_0/n63 ), .A1(\add_x_19_0/n67 ), 
        .B0(\add_x_19_0/n64 ), .Y(\add_x_19_0/n62 ) );
  AOI21X1TS \add_x_19_0/U99  ( .A0(\add_x_19_0/n95 ), .A1(\add_x_19_0/n104 ), 
        .B0(\add_x_19_0/n96 ), .Y(\add_x_19_0/n94 ) );
  OAI21X1TS \add_x_19_0/U101  ( .A0(\add_x_19_0/n97 ), .A1(\add_x_19_0/n101 ), 
        .B0(\add_x_19_0/n98 ), .Y(\add_x_19_0/n96 ) );
  OAI21X1TS \add_x_19_0/U115  ( .A0(\add_x_19_0/n105 ), .A1(\add_x_19_0/n111 ), 
        .B0(\add_x_19_0/n106 ), .Y(\add_x_19_0/n104 ) );
  NOR2X1TS \add_x_19_0/U48  ( .A(\add_x_19_0/n66 ), .B(\add_x_19_0/n63 ), .Y(
        \add_x_19_0/n61 ) );
  NOR2X1TS \add_x_19_0/U69  ( .A(\add_x_19_0/n81 ), .B(\add_x_19_0/n78 ), .Y(
        \add_x_19_0/n76 ) );
  NOR2X1TS \add_x_19_0/U100  ( .A(\add_x_19_0/n100 ), .B(\add_x_19_0/n97 ), 
        .Y(\add_x_19_0/n95 ) );
  NOR2X1TS \add_x_19_0/U114  ( .A(\add_x_19_0/n110 ), .B(\add_x_19_0/n105 ), 
        .Y(\add_x_19_0/n103 ) );
  AOI21X1TS \add_x_19_0/U165  ( .A0(\add_x_19_0/n137 ), .A1(\add_x_19_0/n150 ), 
        .B0(\add_x_19_0/n138 ), .Y(\add_x_19_0/n136 ) );
  OAI21X1TS \add_x_19_0/U167  ( .A0(\add_x_19_0/n139 ), .A1(\add_x_19_0/n145 ), 
        .B0(\add_x_19_0/n140 ), .Y(\add_x_19_0/n138 ) );
  OAI21X1TS \add_x_19_0/U185  ( .A0(\add_x_19_0/n151 ), .A1(\add_x_19_0/n155 ), 
        .B0(\add_x_19_0/n152 ), .Y(\add_x_19_0/n150 ) );
  NOR2X1TS \add_x_19_0/U149  ( .A(\add_x_19_0/n131 ), .B(\add_x_19_0/n128 ), 
        .Y(\add_x_19_0/n126 ) );
  NOR2X1TS \add_x_19_0/U166  ( .A(\add_x_19_0/n144 ), .B(\add_x_19_0/n139 ), 
        .Y(\add_x_19_0/n137 ) );
  NOR2X1TS \add_x_19_0/U170  ( .A(\addr_calc/fft_read_calc/count[11] ), .B(
        n2406), .Y(\add_x_19_0/n139 ) );
  NOR2X1TS \add_x_19_0/U184  ( .A(\add_x_19_0/n154 ), .B(\add_x_19_0/n151 ), 
        .Y(\add_x_19_0/n149 ) );
  OAI21X1TS \add_x_19_0/U216  ( .A0(\add_x_19_0/n170 ), .A1(\add_x_19_0/n176 ), 
        .B0(\add_x_19_0/n171 ), .Y(\add_x_19_0/n169 ) );
  NOR2X1TS \add_x_19_0/U215  ( .A(\add_x_19_0/n175 ), .B(\add_x_19_0/n170 ), 
        .Y(\add_x_19_0/n168 ) );
  NOR2X1TS \add_x_19_0/U249  ( .A(\addr_calc/fft_read_calc/count[1] ), .B(
        n2454), .Y(\add_x_19_0/n188 ) );
  XOR2X1TS \add_x_19_0/U112  ( .A(\add_x_19_0/n107 ), .B(\add_x_19_0/n15 ), 
        .Y(\addr_calc/fft_read_addr[17] ) );
  NAND2X1TS \add_x_19_0/U11  ( .A(\addr_calc/fft_read_calc/count[30] ), .B(
        n2457), .Y(\add_x_19_0/n37 ) );
  NAND2X1TS \add_x_19_0/U19  ( .A(n1863), .B(n2389), .Y(\add_x_19_0/n42 ) );
  NAND2X1TS \add_x_19_0/U29  ( .A(n2559), .B(n2385), .Y(\add_x_19_0/n49 ) );
  NAND2X1TS \add_x_19_0/U39  ( .A(n1944), .B(n2500), .Y(\add_x_19_0/n56 ) );
  NAND2X1TS \add_x_19_0/U45  ( .A(\addr_calc/fft_read_calc/count[26] ), .B(
        n2377), .Y(\add_x_19_0/n59 ) );
  NAND2X1TS \add_x_19_0/U53  ( .A(n1947), .B(n2491), .Y(\add_x_19_0/n64 ) );
  NAND2X1TS \add_x_19_0/U59  ( .A(n2038), .B(n2461), .Y(\add_x_19_0/n67 ) );
  NAND2X1TS \add_x_19_0/U74  ( .A(n1950), .B(n2469), .Y(\add_x_19_0/n79 ) );
  NAND2X1TS \add_x_19_0/U80  ( .A(\addr_calc/fft_read_calc/count[22] ), .B(
        n2466), .Y(\add_x_19_0/n82 ) );
  NAND2X1TS \add_x_19_0/U88  ( .A(\addr_calc/fft_read_calc/count[21] ), .B(
        n2448), .Y(\add_x_19_0/n87 ) );
  NAND2X1TS \add_x_19_0/U105  ( .A(n1956), .B(n2488), .Y(\add_x_19_0/n98 ) );
  NAND2X1TS \add_x_19_0/U111  ( .A(\addr_calc/fft_read_calc/count[18] ), .B(
        n2432), .Y(\add_x_19_0/n101 ) );
  NAND2X1TS \add_x_19_0/U119  ( .A(n1960), .B(n2481), .Y(\add_x_19_0/n106 ) );
  NOR2X1TS \add_x_19_0/U52  ( .A(n1947), .B(n2492), .Y(\add_x_19_0/n63 ) );
  NOR2X1TS \add_x_19_0/U58  ( .A(n2038), .B(n2460), .Y(\add_x_19_0/n66 ) );
  NOR2X1TS \add_x_19_0/U79  ( .A(n1665), .B(n2466), .Y(\add_x_19_0/n81 ) );
  NOR2X1TS \add_x_19_0/U87  ( .A(\addr_calc/fft_read_calc/count[21] ), .B(
        n2449), .Y(\add_x_19_0/n86 ) );
  NOR2X1TS \add_x_19_0/U110  ( .A(\addr_calc/fft_read_calc/count[18] ), .B(
        n2432), .Y(\add_x_19_0/n100 ) );
  NOR2X1TS \add_x_19_0/U118  ( .A(n1960), .B(n2481), .Y(\add_x_19_0/n105 ) );
  NAND2X1TS \add_x_19_0/U140  ( .A(n1689), .B(n2477), .Y(\add_x_19_0/n121 ) );
  NAND2X1TS \add_x_19_0/U146  ( .A(n2043), .B(n2425), .Y(\add_x_19_0/n124 ) );
  NAND2X1TS \add_x_19_0/U154  ( .A(n1967), .B(n2416), .Y(\add_x_19_0/n129 ) );
  NAND2X1TS \add_x_19_0/U179  ( .A(n2413), .B(
        \addr_calc/fft_read_calc/count[10] ), .Y(\add_x_19_0/n145 ) );
  NAND2X1TS \add_x_19_0/U189  ( .A(\addr_calc/fft_read_calc/count[9] ), .B(
        n2496), .Y(\add_x_19_0/n152 ) );
  NAND2X1TS \add_x_19_0/U195  ( .A(\addr_calc/fft_read_calc/count[8] ), .B(
        n2473), .Y(\add_x_19_0/n155 ) );
  NOR2X1TS \add_x_19_0/U159  ( .A(n2046), .B(n2409), .Y(\add_x_19_0/n131 ) );
  NOR2X1TS \add_x_19_0/U178  ( .A(\addr_calc/fft_read_calc/count[10] ), .B(
        n2413), .Y(\add_x_19_0/n144 ) );
  NOR2X1TS \add_x_19_0/U188  ( .A(\addr_calc/fft_read_calc/count[9] ), .B(
        n2495), .Y(\add_x_19_0/n151 ) );
  NOR2X1TS \add_x_19_0/U194  ( .A(\addr_calc/fft_read_calc/count[8] ), .B(
        n2473), .Y(\add_x_19_0/n154 ) );
  NAND2X1TS \add_x_19_0/U206  ( .A(n1666), .B(n2422), .Y(\add_x_19_0/n163 ) );
  NAND2X1TS \add_x_19_0/U212  ( .A(\addr_calc/fft_read_calc/count[6] ), .B(
        n2430), .Y(\add_x_19_0/n166 ) );
  NAND2X1TS \add_x_19_0/U228  ( .A(\addr_calc/fft_read_calc/count[4] ), .B(
        n2397), .Y(\add_x_19_0/n176 ) );
  NAND2X1TS \add_x_19_0/U237  ( .A(\addr_calc/fft_read_calc/count[3] ), .B(
        n2436), .Y(\add_x_19_0/n182 ) );
  NAND2X1TS \add_x_19_0/U243  ( .A(\addr_calc/fft_read_calc/count[2] ), .B(
        n2445), .Y(\add_x_19_0/n185 ) );
  NAND2X1TS \add_x_19_0/U250  ( .A(\addr_calc/fft_read_calc/count[1] ), .B(
        n2453), .Y(\add_x_19_0/n189 ) );
  NOR2X1TS \add_x_19_0/U242  ( .A(\addr_calc/fft_read_calc/count[2] ), .B(
        n2445), .Y(\add_x_19_0/n184 ) );
  XNOR2X1TS \add_x_19_0/U221  ( .A(\add_x_19_0/n177 ), .B(\add_x_19_0/n28 ), 
        .Y(\addr_calc/fft_read_addr[4] ) );
  NAND2X1TS \add_x_19_0/U225  ( .A(\add_x_19_0/n219 ), .B(\add_x_19_0/n176 ), 
        .Y(\add_x_19_0/n28 ) );
  NAND2X1TS \add_x_19_0/U192  ( .A(\add_x_19_0/n215 ), .B(\add_x_19_0/n155 ), 
        .Y(\add_x_19_0/n24 ) );
  XNOR2X1TS \add_x_19_0/U172  ( .A(\add_x_19_0/n146 ), .B(\add_x_19_0/n22 ), 
        .Y(\addr_calc/fft_read_addr[10] ) );
  NAND2X1TS \add_x_19_0/U176  ( .A(\add_x_19_0/n213 ), .B(\add_x_19_0/n145 ), 
        .Y(\add_x_19_0/n22 ) );
  XNOR2X1TS \add_x_19_0/U147  ( .A(\add_x_19_0/n130 ), .B(\add_x_19_0/n19 ), 
        .Y(\addr_calc/fft_read_addr[13] ) );
  NAND2X1TS \add_x_19_0/U151  ( .A(\add_x_19_0/n210 ), .B(\add_x_19_0/n129 ), 
        .Y(\add_x_19_0/n19 ) );
  XNOR2X1TS \add_x_19_0/U128  ( .A(\add_x_19_0/n122 ), .B(\add_x_19_0/n17 ), 
        .Y(\addr_calc/fft_read_addr[15] ) );
  NAND2X1TS \add_x_19_0/U137  ( .A(\add_x_19_0/n208 ), .B(\add_x_19_0/n121 ), 
        .Y(\add_x_19_0/n17 ) );
  NAND2X1TS \add_x_19_0/U116  ( .A(\add_x_19_0/n206 ), .B(\add_x_19_0/n106 ), 
        .Y(\add_x_19_0/n15 ) );
  XNOR2X1TS \add_x_19_0/U95  ( .A(\add_x_19_0/n99 ), .B(\add_x_19_0/n13 ), .Y(
        \addr_calc/fft_read_addr[19] ) );
  NAND2X1TS \add_x_19_0/U102  ( .A(\add_x_19_0/n204 ), .B(\add_x_19_0/n98 ), 
        .Y(\add_x_19_0/n13 ) );
  XNOR2X1TS \add_x_19_0/U81  ( .A(\add_x_19_0/n88 ), .B(\add_x_19_0/n11 ), .Y(
        \addr_calc/fft_read_addr[21] ) );
  NAND2X1TS \add_x_19_0/U85  ( .A(\add_x_19_0/n202 ), .B(\add_x_19_0/n87 ), 
        .Y(\add_x_19_0/n11 ) );
  NAND2X1TS \add_x_19_0/U26  ( .A(\add_x_19_0/n195 ), .B(\add_x_19_0/n49 ), 
        .Y(\add_x_19_0/n4 ) );
  XNOR2X1TS \add_x_19_0/U46  ( .A(\add_x_19_0/n65 ), .B(\add_x_19_0/n7 ), .Y(
        \addr_calc/fft_read_addr[25] ) );
  NAND2X1TS \add_x_19_0/U50  ( .A(\add_x_19_0/n198 ), .B(\add_x_19_0/n64 ), 
        .Y(\add_x_19_0/n7 ) );
  NAND2X1TS \add_x_19_0/U2  ( .A(n2627), .B(\add_x_19_0/n34 ), .Y(
        \add_x_19_0/n1 ) );
  NAND2X1TS \add_x_19_0/U22  ( .A(\add_x_19_0/n72 ), .B(\add_x_19_0/n46 ), .Y(
        \add_x_19_0/n44 ) );
  NAND2X1TS \add_x_19_0/U32  ( .A(\add_x_19_0/n61 ), .B(\add_x_19_0/n53 ), .Y(
        \add_x_19_0/n51 ) );
  NAND2X1TS \add_x_19_0/U98  ( .A(\add_x_19_0/n103 ), .B(\add_x_19_0/n95 ), 
        .Y(\add_x_19_0/n93 ) );
  NAND2X1TS \add_x_19_0/U171  ( .A(\addr_calc/fft_read_calc/count[11] ), .B(
        n2406), .Y(\add_x_19_0/n140 ) );
  NAND2X1TS \add_x_19_0/U164  ( .A(\add_x_19_0/n149 ), .B(\add_x_19_0/n137 ), 
        .Y(\add_x_19_0/n135 ) );
  NAND2X1TS \add_x_19_0/U220  ( .A(\addr_calc/fft_read_calc/count[5] ), .B(
        n2485), .Y(\add_x_19_0/n171 ) );
  NOR2X2TS \DP_OP_159_297_3515/U1098  ( .A(\DP_OP_159_297_3515/n1063 ), .B(
        \DP_OP_159_297_3515/n1052 ), .Y(\DP_OP_159_297_3515/n1051 ) );
  NAND2X1TS \DP_OP_159_297_3515/U964  ( .A(n1531), .B(n1491), .Y(
        \DP_OP_159_297_3515/n959 ) );
  NOR2XLTS \DP_OP_159_297_3515/U1050  ( .A(\DP_OP_159_297_3515/n1026 ), .B(
        \DP_OP_159_297_3515/n873 ), .Y(\DP_OP_159_297_3515/n1018 ) );
  NAND2X2TS \DP_OP_159_297_3515/U990  ( .A(n1789), .B(n2369), .Y(
        \DP_OP_159_297_3515/n976 ) );
  NOR2X1TS \DP_OP_159_297_3515/U798  ( .A(\DP_OP_159_297_3515/n768 ), .B(
        \DP_OP_159_297_3515/n766 ), .Y(\DP_OP_159_297_3515/n764 ) );
  NOR2X1TS \DP_OP_159_297_3515/U810  ( .A(\DP_OP_159_297_3515/n776 ), .B(
        \DP_OP_159_297_3515/n778 ), .Y(\DP_OP_159_297_3515/n774 ) );
  NOR2X1TS \DP_OP_159_297_3515/U757  ( .A(\DP_OP_159_297_3515/n730 ), .B(
        \DP_OP_159_297_3515/n737 ), .Y(\DP_OP_159_297_3515/n728 ) );
  NOR2X1TS \DP_OP_159_297_3515/U1030  ( .A(\DP_OP_159_297_3515/n1012 ), .B(
        \DP_OP_159_297_3515/n871 ), .Y(\DP_OP_159_297_3515/n1004 ) );
  NOR2X1TS \DP_OP_159_297_3515/U1020  ( .A(\DP_OP_159_297_3515/n1012 ), .B(
        \DP_OP_159_297_3515/n998 ), .Y(\DP_OP_159_297_3515/n997 ) );
  NOR2X1TS \DP_OP_159_297_3515/U971  ( .A(\DP_OP_159_297_3515/n971 ), .B(
        \DP_OP_159_297_3515/n964 ), .Y(\DP_OP_159_297_3515/n963 ) );
  NOR2X1TS \DP_OP_159_297_3515/U861  ( .A(n2551), .B(\DP_OP_159_297_3515/n887 ), .Y(\DP_OP_159_297_3515/n886 ) );
  NOR2X1TS \DP_OP_159_297_3515/U871  ( .A(\DP_OP_159_297_3515/n852 ), .B(
        \DP_OP_159_297_3515/n894 ), .Y(\DP_OP_159_297_3515/n893 ) );
  NOR2X1TS \DP_OP_159_297_3515/U931  ( .A(\DP_OP_159_297_3515/n957 ), .B(
        \DP_OP_159_297_3515/n936 ), .Y(\DP_OP_159_297_3515/n935 ) );
  NOR2X1TS \DP_OP_159_297_3515/U951  ( .A(\DP_OP_159_297_3515/n957 ), .B(
        \DP_OP_159_297_3515/n950 ), .Y(\DP_OP_159_297_3515/n949 ) );
  NOR2X1TS \DP_OP_159_297_3515/U891  ( .A(n2551), .B(\DP_OP_159_297_3515/n908 ), .Y(\DP_OP_159_297_3515/n907 ) );
  NOR2X1TS \DP_OP_159_297_3515/U901  ( .A(\DP_OP_159_297_3515/n852 ), .B(
        \DP_OP_159_297_3515/n915 ), .Y(\DP_OP_159_297_3515/n914 ) );
  NAND2X1TS \DP_OP_159_297_3515/U791  ( .A(\DP_OP_159_297_3515/n764 ), .B(
        n2606), .Y(\DP_OP_159_297_3515/n758 ) );
  XNOR2X1TS \DP_OP_159_297_3515/U800  ( .A(n2611), .B(
        \addr_calc/iir_write_calc/count[3] ), .Y(\DP_OP_159_297_3515/n766 ) );
  NAND2X1TS \DP_OP_159_297_3515/U803  ( .A(\DP_OP_159_297_3515/n774 ), .B(
        n2604), .Y(\DP_OP_159_297_3515/n768 ) );
  XNOR2X1TS \DP_OP_159_297_3515/U812  ( .A(n2374), .B(
        \addr_calc/iir_write_calc/count[1] ), .Y(\DP_OP_159_297_3515/n776 ) );
  NAND2X1TS \DP_OP_159_297_3515/U773  ( .A(n2605), .B(n2626), .Y(
        \DP_OP_159_297_3515/n742 ) );
  XNOR2X1TS \DP_OP_159_297_3515/U767  ( .A(n2609), .B(
        \addr_calc/iir_write_calc/count[7] ), .Y(\DP_OP_159_297_3515/n737 ) );
  NAND2X1TS \DP_OP_159_297_3515/U1088  ( .A(\DP_OP_159_297_3515/n1051 ), .B(
        n2362), .Y(\DP_OP_159_297_3515/n1044 ) );
  NAND2X1TS \DP_OP_159_297_3515/U1011  ( .A(\DP_OP_159_297_3515/n999 ), .B(
        n1521), .Y(\DP_OP_159_297_3515/n991 ) );
  NAND2X1TS \DP_OP_159_297_3515/U860  ( .A(n1790), .B(
        \DP_OP_159_297_3515/n886 ), .Y(\DP_OP_159_297_3515/n885 ) );
  NAND2X1TS \DP_OP_159_297_3515/U862  ( .A(\DP_OP_159_297_3515/n902 ), .B(
        n2603), .Y(\DP_OP_159_297_3515/n887 ) );
  NAND2X1TS \DP_OP_159_297_3515/U872  ( .A(\DP_OP_159_297_3515/n902 ), .B(
        n2342), .Y(\DP_OP_159_297_3515/n894 ) );
  NAND2X1TS \DP_OP_159_297_3515/U932  ( .A(\DP_OP_159_297_3515/n944 ), .B(
        n2344), .Y(\DP_OP_159_297_3515/n936 ) );
  NAND2X1TS \DP_OP_159_297_3515/U892  ( .A(\DP_OP_159_297_3515/n916 ), .B(
        n1562), .Y(\DP_OP_159_297_3515/n908 ) );
  NAND2X1TS \DP_OP_159_297_3515/U924  ( .A(n1518), .B(n1815), .Y(
        \DP_OP_159_297_3515/n931 ) );
  NOR2X2TS \DP_OP_158_296_6262/U305  ( .A(\DP_OP_158_296_6262/n282 ), .B(
        \DP_OP_158_296_6262/n318 ), .Y(\DP_OP_158_296_6262/n280 ) );
  NOR2X1TS \DP_OP_158_296_6262/U379  ( .A(\DP_OP_158_296_6262/n349 ), .B(
        \DP_OP_158_296_6262/n365 ), .Y(\DP_OP_158_296_6262/n347 ) );
  NOR2X1TS \DP_OP_158_296_6262/U406  ( .A(\DP_OP_158_296_6262/n373 ), .B(
        \DP_OP_158_296_6262/n375 ), .Y(\DP_OP_158_296_6262/n371 ) );
  NOR2X1TS \DP_OP_158_296_6262/U309  ( .A(\DP_OP_158_296_6262/n297 ), .B(
        \DP_OP_158_296_6262/n286 ), .Y(\DP_OP_158_296_6262/n284 ) );
  NOR2X1TS \DP_OP_158_296_6262/U1803  ( .A(\DP_OP_158_296_6262/n1792 ), .B(
        \DP_OP_158_296_6262/n1829 ), .Y(\DP_OP_158_296_6262/n1828 ) );
  NAND2X1TS \DP_OP_158_296_6262/U399  ( .A(\DP_OP_158_296_6262/n371 ), .B(
        n2590), .Y(\DP_OP_158_296_6262/n365 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U408  ( .A(n2597), .B(n1910), .Y(
        \DP_OP_158_296_6262/n373 ) );
  NAND2X1TS \DP_OP_158_296_6262/U381  ( .A(n2592), .B(n2600), .Y(
        \DP_OP_158_296_6262/n349 ) );
  NAND2X1TS \DP_OP_158_296_6262/U359  ( .A(n2601), .B(n2591), .Y(
        \DP_OP_158_296_6262/n329 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U351  ( .A(n1651), .B(n1480), .Y(
        \DP_OP_158_296_6262/n322 ) );
  NAND2X1TS \DP_OP_158_296_6262/U307  ( .A(\DP_OP_158_296_6262/n284 ), .B(
        \DP_OP_158_296_6262/n304 ), .Y(\DP_OP_158_296_6262/n282 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U343  ( .A(n2598), .B(n1997), .Y(
        \DP_OP_158_296_6262/n315 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U333  ( .A(n1469), .B(n1900), .Y(
        \DP_OP_158_296_6262/n306 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U311  ( .A(n1660), .B(n1895), .Y(
        \DP_OP_158_296_6262/n286 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U263  ( .A(n1658), .B(n1890), .Y(
        \DP_OP_158_296_6262/n242 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U277  ( .A(n1657), .B(n1690), .Y(
        \DP_OP_158_296_6262/n255 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U289  ( .A(n1659), .B(n1893), .Y(
        \DP_OP_158_296_6262/n266 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U250  ( .A(n2594), .B(n1888), .Y(
        \DP_OP_158_296_6262/n230 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U10  ( .A(n1778), .B(
        \addr_calc/fir_read_calc/count[31] ), .Y(\DP_OP_158_296_6262/n5 ) );
  NAND2X1TS \DP_OP_158_296_6262/U2032  ( .A(\DP_OP_158_296_6262/n2010 ), .B(
        \DP_OP_159_297_3515/n880 ), .Y(\DP_OP_158_296_6262/n2004 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1981  ( .A(n1138), .B(
        \DP_OP_158_296_6262/n1966 ), .Y(\DP_OP_158_296_6262/n1965 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1945  ( .A(\DP_OP_158_296_6262/n1938 ), .B(
        \DP_OP_158_296_6262/n1959 ), .Y(\DP_OP_158_296_6262/n1937 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1963  ( .A(\DP_OP_158_296_6262/n1959 ), .B(
        \DP_OP_158_296_6262/n1952 ), .Y(\DP_OP_158_296_6262/n1951 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1910  ( .A(\DP_OP_158_296_6262/n1918 ), .B(
        \DP_OP_158_296_6262/n1911 ), .Y(\DP_OP_158_296_6262/n1910 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1802  ( .A(\DP_OP_158_296_6262/n1791 ), .B(
        \DP_OP_158_296_6262/n1828 ), .Y(\DP_OP_158_296_6262/n1827 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1838  ( .A(\DP_OP_158_296_6262/n1855 ), .B(
        n1783), .Y(\DP_OP_158_296_6262/n1854 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1892  ( .A(\DP_OP_158_296_6262/n1904 ), .B(
        \DP_OP_158_296_6262/n1897 ), .Y(\DP_OP_158_296_6262/n1896 ) );
  NOR2X1TS \add_x_22_4/U101  ( .A(\add_x_22_4/n85 ), .B(\add_x_22_4/n84 ), .Y(
        \add_x_22_4/n81 ) );
  NOR2X1TS \add_x_22_4/U127  ( .A(\add_x_22_4/n110 ), .B(\add_x_22_4/n103 ), 
        .Y(\add_x_22_4/n102 ) );
  NOR2X1TS \add_x_22_4/U132  ( .A(\add_x_22_4/n110 ), .B(\add_x_22_4/n109 ), 
        .Y(\add_x_22_4/n106 ) );
  NOR2X1TS \add_x_22_4/U85  ( .A(\add_x_22_4/n76 ), .B(\add_x_22_4/n69 ), .Y(
        \add_x_22_4/n68 ) );
  NOR2X1TS \add_x_22_4/U63  ( .A(\add_x_22_4/n58 ), .B(\add_x_22_4/n51 ), .Y(
        \add_x_22_4/n50 ) );
  NOR2X1TS \add_x_22_4/U21  ( .A(\add_x_22_4/n24 ), .B(\add_x_22_4/n17 ), .Y(
        \add_x_22_4/n16 ) );
  NOR2X1TS \add_x_22_4/U12  ( .A(\add_x_22_4/n17 ), .B(\add_x_22_4/n10 ), .Y(
        \add_x_22_4/n9 ) );
  NOR2X1TS \add_x_22_4/U34  ( .A(\add_x_22_4/n35 ), .B(\add_x_22_4/n28 ), .Y(
        \add_x_22_4/n27 ) );
  NOR2X1TS \add_x_22_4/U68  ( .A(\add_x_22_4/n58 ), .B(\add_x_22_4/n57 ), .Y(
        \add_x_22_4/n54 ) );
  NOR2X1TS \add_x_22_4/U43  ( .A(\add_x_22_4/n42 ), .B(\add_x_22_4/n35 ), .Y(
        \add_x_22_4/n34 ) );
  NOR2X1TS \add_x_22_4/U54  ( .A(\add_x_22_4/n51 ), .B(\add_x_22_4/n44 ), .Y(
        \add_x_22_4/n43 ) );
  NOR2X1TS \add_x_22_4/U138  ( .A(\add_x_22_4/n112 ), .B(\add_x_22_4/n119 ), 
        .Y(\add_x_22_4/n111 ) );
  NOR2X1TS \add_x_22_4/U96  ( .A(\add_x_22_4/n87 ), .B(\add_x_22_4/n78 ), .Y(
        \add_x_22_4/n77 ) );
  XNOR2X1TS \add_x_22_4/U142  ( .A(\add_x_22_4/n118 ), .B(\add_x_22_4/n117 ), 
        .Y(\addr_calc/iir_read_calc/counter/N45 ) );
  XNOR2X1TS \add_x_22_4/U146  ( .A(\add_x_22_4/n121 ), .B(n2580), .Y(
        \addr_calc/iir_read_calc/counter/N44 ) );
  XNOR2X1TS \add_x_22_4/U80  ( .A(\add_x_22_4/n68 ), .B(\add_x_22_4/n67 ), .Y(
        \addr_calc/iir_read_calc/counter/N57 ) );
  NAND2X1TS \add_x_22_4/U143  ( .A(\add_x_22_4/n118 ), .B(n2015), .Y(
        \add_x_22_4/n115 ) );
  XNOR2X1TS \add_x_22_4/U58  ( .A(\add_x_22_4/n50 ), .B(n2024), .Y(
        \addr_calc/iir_read_calc/counter/N61 ) );
  XNOR2X1TS \add_x_22_4/U47  ( .A(\add_x_22_4/n41 ), .B(n2027), .Y(
        \addr_calc/iir_read_calc/counter/N63 ) );
  XNOR2X1TS \add_x_22_4/U89  ( .A(\add_x_22_4/n75 ), .B(\add_x_22_4/n74 ), .Y(
        \addr_calc/iir_read_calc/counter/N55 ) );
  XNOR2X1TS \add_x_22_4/U93  ( .A(\add_x_22_4/n81 ), .B(\add_x_22_4/n80 ), .Y(
        \addr_calc/iir_read_calc/counter/N54 ) );
  NAND2X1TS \add_x_22_4/U123  ( .A(\add_x_22_4/n102 ), .B(n2018), .Y(
        \add_x_22_4/n99 ) );
  XNOR2X1TS \add_x_22_4/U126  ( .A(\add_x_22_4/n106 ), .B(\add_x_22_4/n105 ), 
        .Y(\addr_calc/iir_read_calc/counter/N48 ) );
  XNOR2X1TS \add_x_22_4/U111  ( .A(\add_x_22_4/n93 ), .B(\add_x_22_4/n92 ), 
        .Y(\addr_calc/iir_read_calc/counter/N51 ) );
  NAND2X1TS \add_x_22_4/U81  ( .A(\add_x_22_4/n68 ), .B(n1784), .Y(
        \add_x_22_4/n65 ) );
  NAND2X1TS \add_x_22_4/U95  ( .A(\add_x_22_4/n93 ), .B(\add_x_22_4/n77 ), .Y(
        \add_x_22_4/n76 ) );
  NAND2X1TS \add_x_22_4/U11  ( .A(\add_x_22_4/n23 ), .B(\add_x_22_4/n9 ), .Y(
        \add_x_22_4/n8 ) );
  NAND2X1TS \add_x_22_4/U59  ( .A(\add_x_22_4/n50 ), .B(
        \addr_calc/iir_read_calc/count[18] ), .Y(\add_x_22_4/n47 ) );
  NAND2X1TS \add_x_22_4/U26  ( .A(\add_x_22_4/n23 ), .B(n2034), .Y(
        \add_x_22_4/n20 ) );
  XNOR2X1TS \add_x_22_4/U25  ( .A(\add_x_22_4/n23 ), .B(n2033), .Y(
        \addr_calc/iir_read_calc/counter/N67 ) );
  ADDHXLTS \add_x_22_4/U2  ( .A(\addr_calc/iir_read_calc/count[30] ), .B(
        \add_x_22_4/n2 ), .CO(\add_x_22_4/n1 ), .S(
        \addr_calc/iir_read_calc/counter/N73 ) );
  NAND2X1TS \add_x_22_4/U13  ( .A(n2576), .B(n1929), .Y(\add_x_22_4/n10 ) );
  NAND2X1TS \add_x_22_4/U22  ( .A(\addr_calc/iir_read_calc/count[24] ), .B(
        n1926), .Y(\add_x_22_4/n17 ) );
  NAND2X1TS \add_x_22_4/U33  ( .A(\add_x_22_4/n43 ), .B(\add_x_22_4/n27 ), .Y(
        \add_x_22_4/n26 ) );
  NAND2X1TS \add_x_22_4/U35  ( .A(n2031), .B(n2565), .Y(\add_x_22_4/n28 ) );
  XNOR2X1TS \add_x_22_4/U62  ( .A(\add_x_22_4/n54 ), .B(n1919), .Y(
        \addr_calc/iir_read_calc/counter/N60 ) );
  NAND2X1TS \add_x_22_4/U44  ( .A(n2028), .B(n1687), .Y(\add_x_22_4/n35 ) );
  NAND2X1TS \add_x_22_4/U53  ( .A(\add_x_22_4/n59 ), .B(\add_x_22_4/n43 ), .Y(
        \add_x_22_4/n42 ) );
  NAND2X1TS \add_x_22_4/U55  ( .A(n2025), .B(
        \addr_calc/iir_read_calc/count[19] ), .Y(\add_x_22_4/n44 ) );
  NAND2X1TS \add_x_22_4/U64  ( .A(\addr_calc/iir_read_calc/count[16] ), .B(
        n1920), .Y(\add_x_22_4/n51 ) );
  NAND2X1TS \add_x_22_4/U148  ( .A(n1898), .B(
        \addr_calc/iir_read_calc/count[0] ), .Y(\add_x_22_4/n119 ) );
  NAND2X1TS \add_x_22_4/U139  ( .A(n2015), .B(
        \addr_calc/iir_read_calc/count[3] ), .Y(\add_x_22_4/n112 ) );
  NAND2X1TS \add_x_22_4/U128  ( .A(\addr_calc/iir_read_calc/count[4] ), .B(
        \addr_calc/iir_read_calc/count[5] ), .Y(\add_x_22_4/n103 ) );
  NAND2X1TS \add_x_22_4/U86  ( .A(\addr_calc/iir_read_calc/count[12] ), .B(
        \addr_calc/iir_read_calc/count[13] ), .Y(\add_x_22_4/n69 ) );
  NAND2X1TS \add_x_22_4/U97  ( .A(n1909), .B(n1911), .Y(\add_x_22_4/n78 ) );
  NAND2X1TS \add_x_22_4/U108  ( .A(\addr_calc/iir_read_calc/count[8] ), .B(
        n1685), .Y(\add_x_22_4/n87 ) );
  XOR2X1TS \add_x_22_4/U136  ( .A(\add_x_22_4/n115 ), .B(n1901), .Y(
        \addr_calc/iir_read_calc/counter/N46 ) );
  XOR2X1TS \add_x_22_4/U115  ( .A(\add_x_22_4/n99 ), .B(\add_x_22_4/n98 ), .Y(
        \addr_calc/iir_read_calc/counter/N50 ) );
  XOR2X1TS \add_x_22_4/U105  ( .A(\add_x_22_4/n90 ), .B(n1907), .Y(
        \addr_calc/iir_read_calc/counter/N52 ) );
  XOR2X1TS \add_x_22_4/U100  ( .A(\add_x_22_4/n85 ), .B(\add_x_22_4/n84 ), .Y(
        \addr_calc/iir_read_calc/counter/N53 ) );
  XOR2X1TS \add_x_22_4/U72  ( .A(\add_x_22_4/n65 ), .B(\add_x_22_4/n64 ), .Y(
        \addr_calc/iir_read_calc/counter/N58 ) );
  XOR2X1TS \add_x_22_4/U67  ( .A(\add_x_22_4/n58 ), .B(\add_x_22_4/n57 ), .Y(
        \addr_calc/iir_read_calc/counter/N59 ) );
  XOR2X1TS \add_x_22_4/U51  ( .A(\add_x_22_4/n47 ), .B(\add_x_22_4/n46 ), .Y(
        \addr_calc/iir_read_calc/counter/N62 ) );
  XOR2X1TS \add_x_22_4/U20  ( .A(\add_x_22_4/n20 ), .B(n1925), .Y(
        \addr_calc/iir_read_calc/counter/N68 ) );
  XOR2X1TS \add_x_22_4/U4  ( .A(\add_x_22_4/n8 ), .B(\add_x_22_4/n7 ), .Y(
        \addr_calc/iir_read_calc/counter/N71 ) );
  XOR2X1TS \add_x_22_4/U1  ( .A(\add_x_22_4/n1 ), .B(
        \addr_calc/iir_read_calc/count[31] ), .Y(
        \addr_calc/iir_read_calc/counter/N74 ) );
  NOR2X1TS \add_x_22_1/U127  ( .A(\add_x_22_1/n110 ), .B(\add_x_22_1/n103 ), 
        .Y(\add_x_22_1/n102 ) );
  NOR2X1TS \add_x_22_1/U85  ( .A(\add_x_22_1/n76 ), .B(\add_x_22_1/n69 ), .Y(
        \add_x_22_1/n68 ) );
  NOR2X1TS \add_x_22_1/U63  ( .A(\add_x_22_1/n58 ), .B(\add_x_22_1/n51 ), .Y(
        \add_x_22_1/n50 ) );
  NOR2X1TS \add_x_22_1/U68  ( .A(\add_x_22_1/n58 ), .B(\add_x_22_1/n57 ), .Y(
        \add_x_22_1/n54 ) );
  NOR2X1TS \add_x_22_1/U43  ( .A(\add_x_22_1/n42 ), .B(\add_x_22_1/n35 ), .Y(
        \add_x_22_1/n34 ) );
  NOR2X1TS \add_x_22_1/U21  ( .A(\add_x_22_1/n24 ), .B(\add_x_22_1/n17 ), .Y(
        \add_x_22_1/n16 ) );
  NOR2X1TS \add_x_22_1/U6  ( .A(\add_x_22_1/n26 ), .B(\add_x_22_1/n5 ), .Y(
        \add_x_22_1/n4 ) );
  NOR2X1TS \add_x_22_1/U12  ( .A(\add_x_22_1/n17 ), .B(\add_x_22_1/n10 ), .Y(
        \add_x_22_1/n9 ) );
  NOR2X1TS \add_x_22_1/U34  ( .A(\add_x_22_1/n35 ), .B(\add_x_22_1/n28 ), .Y(
        \add_x_22_1/n27 ) );
  NOR2X1TS \add_x_22_1/U54  ( .A(\add_x_22_1/n51 ), .B(\add_x_22_1/n44 ), .Y(
        \add_x_22_1/n43 ) );
  NOR2X1TS \add_x_22_1/U138  ( .A(\add_x_22_1/n112 ), .B(\add_x_22_1/n119 ), 
        .Y(\add_x_22_1/n111 ) );
  NOR2X1TS \add_x_22_1/U118  ( .A(\add_x_22_1/n103 ), .B(\add_x_22_1/n96 ), 
        .Y(\add_x_22_1/n95 ) );
  NOR2X1TS \add_x_22_1/U96  ( .A(\add_x_22_1/n87 ), .B(\add_x_22_1/n78 ), .Y(
        \add_x_22_1/n77 ) );
  NAND2X1TS \add_x_22_1/U90  ( .A(\add_x_22_1/n75 ), .B(n2023), .Y(
        \add_x_22_1/n72 ) );
  XNOR2X1TS \add_x_22_1/U89  ( .A(\add_x_22_1/n75 ), .B(\add_x_22_1/n74 ), .Y(
        \addr_calc/fft_write_calc/counter/N55 ) );
  NAND2X1TS \add_x_22_1/U123  ( .A(\add_x_22_1/n102 ), .B(n2030), .Y(
        \add_x_22_1/n99 ) );
  XNOR2X1TS \add_x_22_1/U111  ( .A(\add_x_22_1/n93 ), .B(\add_x_22_1/n92 ), 
        .Y(\addr_calc/fft_write_calc/counter/N51 ) );
  XNOR2X1TS \add_x_22_1/U80  ( .A(\add_x_22_1/n68 ), .B(\add_x_22_1/n67 ), .Y(
        \addr_calc/fft_write_calc/counter/N57 ) );
  NAND2X1TS \add_x_22_1/U143  ( .A(\add_x_22_1/n118 ), .B(n2032), .Y(
        \add_x_22_1/n115 ) );
  NAND2X1TS \add_x_22_1/U95  ( .A(\add_x_22_1/n93 ), .B(\add_x_22_1/n77 ), .Y(
        \add_x_22_1/n76 ) );
  NAND2X1TS \add_x_22_1/U48  ( .A(\add_x_22_1/n41 ), .B(
        \addr_calc/fft_write_calc/count[20] ), .Y(\add_x_22_1/n38 ) );
  XNOR2X1TS \add_x_22_1/U62  ( .A(\add_x_22_1/n54 ), .B(\add_x_22_1/n53 ), .Y(
        \addr_calc/fft_write_calc/counter/N60 ) );
  NAND2X1TS \add_x_22_1/U53  ( .A(\add_x_22_1/n59 ), .B(\add_x_22_1/n43 ), .Y(
        \add_x_22_1/n42 ) );
  NAND2X1TS \add_x_22_1/U26  ( .A(\add_x_22_1/n23 ), .B(
        \addr_calc/fft_write_calc/count[24] ), .Y(\add_x_22_1/n20 ) );
  NAND2X1TS \add_x_22_1/U11  ( .A(\add_x_22_1/n23 ), .B(\add_x_22_1/n9 ), .Y(
        \add_x_22_1/n8 ) );
  ADDHXLTS \add_x_22_1/U2  ( .A(\addr_calc/fft_write_calc/count[30] ), .B(
        \add_x_22_1/n2 ), .CO(\add_x_22_1/n1 ), .S(
        \addr_calc/fft_write_calc/counter/N73 ) );
  NAND2X1TS \add_x_22_1/U22  ( .A(n2011), .B(
        \addr_calc/fft_write_calc/count[25] ), .Y(\add_x_22_1/n17 ) );
  NAND2X1TS \add_x_22_1/U33  ( .A(\add_x_22_1/n43 ), .B(\add_x_22_1/n27 ), .Y(
        \add_x_22_1/n26 ) );
  NAND2X1TS \add_x_22_1/U35  ( .A(n2014), .B(n2555), .Y(\add_x_22_1/n28 ) );
  NAND2X1TS \add_x_22_1/U44  ( .A(n2017), .B(
        \addr_calc/fft_write_calc/count[21] ), .Y(\add_x_22_1/n35 ) );
  NAND2X1TS \add_x_22_1/U55  ( .A(n2020), .B(
        \addr_calc/fft_write_calc/count[19] ), .Y(\add_x_22_1/n44 ) );
  NAND2X1TS \add_x_22_1/U64  ( .A(n2567), .B(n1924), .Y(\add_x_22_1/n51 ) );
  NAND2X1TS \add_x_22_1/U117  ( .A(\add_x_22_1/n95 ), .B(\add_x_22_1/n111 ), 
        .Y(\add_x_22_1/n94 ) );
  NAND2X1TS \add_x_22_1/U148  ( .A(\addr_calc/fft_write_calc/count[1] ), .B(
        \addr_calc/fft_write_calc/count[0] ), .Y(\add_x_22_1/n119 ) );
  NAND2X1TS \add_x_22_1/U139  ( .A(\addr_calc/fft_write_calc/count[2] ), .B(
        \addr_calc/fft_write_calc/count[3] ), .Y(\add_x_22_1/n112 ) );
  NAND2X1TS \add_x_22_1/U119  ( .A(\addr_calc/fft_write_calc/count[6] ), .B(
        \addr_calc/fft_write_calc/count[7] ), .Y(\add_x_22_1/n96 ) );
  NAND2X1TS \add_x_22_1/U86  ( .A(\addr_calc/fft_write_calc/count[12] ), .B(
        \addr_calc/fft_write_calc/count[13] ), .Y(\add_x_22_1/n69 ) );
  NAND2X1TS \add_x_22_1/U97  ( .A(\addr_calc/fft_write_calc/count[10] ), .B(
        \addr_calc/fft_write_calc/count[11] ), .Y(\add_x_22_1/n78 ) );
  NAND2X1TS \add_x_22_1/U108  ( .A(\addr_calc/fft_write_calc/count[8] ), .B(
        \addr_calc/fft_write_calc/count[9] ), .Y(\add_x_22_1/n87 ) );
  XOR2X1TS \add_x_22_1/U136  ( .A(\add_x_22_1/n115 ), .B(\add_x_22_1/n114 ), 
        .Y(\addr_calc/fft_write_calc/counter/N46 ) );
  XOR2X1TS \add_x_22_1/U131  ( .A(\add_x_22_1/n110 ), .B(\add_x_22_1/n109 ), 
        .Y(\addr_calc/fft_write_calc/counter/N47 ) );
  XOR2X1TS \add_x_22_1/U115  ( .A(\add_x_22_1/n99 ), .B(\add_x_22_1/n98 ), .Y(
        \addr_calc/fft_write_calc/counter/N50 ) );
  XOR2X1TS \add_x_22_1/U105  ( .A(\add_x_22_1/n90 ), .B(\add_x_22_1/n89 ), .Y(
        \addr_calc/fft_write_calc/counter/N52 ) );
  XOR2X1TS \add_x_22_1/U100  ( .A(\add_x_22_1/n85 ), .B(\add_x_22_1/n84 ), .Y(
        \addr_calc/fft_write_calc/counter/N53 ) );
  XOR2X1TS \add_x_22_1/U84  ( .A(\add_x_22_1/n72 ), .B(\add_x_22_1/n71 ), .Y(
        \addr_calc/fft_write_calc/counter/N56 ) );
  XOR2X1TS \add_x_22_1/U72  ( .A(\add_x_22_1/n65 ), .B(\add_x_22_1/n64 ), .Y(
        \addr_calc/fft_write_calc/counter/N58 ) );
  XOR2X1TS \add_x_22_1/U67  ( .A(\add_x_22_1/n58 ), .B(\add_x_22_1/n57 ), .Y(
        \addr_calc/fft_write_calc/counter/N59 ) );
  XOR2X1TS \add_x_22_1/U51  ( .A(\add_x_22_1/n47 ), .B(n1921), .Y(
        \addr_calc/fft_write_calc/counter/N62 ) );
  XOR2X1TS \add_x_22_1/U42  ( .A(\add_x_22_1/n38 ), .B(n1917), .Y(
        \addr_calc/fft_write_calc/counter/N64 ) );
  XOR2X1TS \add_x_22_1/U29  ( .A(\add_x_22_1/n31 ), .B(\add_x_22_1/n30 ), .Y(
        \addr_calc/fft_write_calc/counter/N66 ) );
  XOR2X1TS \add_x_22_1/U20  ( .A(\add_x_22_1/n20 ), .B(n1914), .Y(
        \addr_calc/fft_write_calc/counter/N68 ) );
  XOR2X1TS \add_x_22_1/U4  ( .A(\add_x_22_1/n8 ), .B(\add_x_22_1/n7 ), .Y(
        \addr_calc/fft_write_calc/counter/N71 ) );
  AHHCINX2TS \add_x_22_1/U3  ( .A(\addr_calc/fft_write_calc/count[29] ), .CIN(
        \add_x_22_1/n3 ), .S(\addr_calc/fft_write_calc/counter/N72 ), .CO(
        \add_x_22_1/n2 ) );
  XOR2X1TS \add_x_22_1/U1  ( .A(\add_x_22_1/n1 ), .B(n1845), .Y(
        \addr_calc/fft_write_calc/counter/N74 ) );
  NOR2X1TS \add_x_22_5/U101  ( .A(\add_x_22_5/n85 ), .B(\add_x_22_5/n84 ), .Y(
        \add_x_22_5/n81 ) );
  NOR2X1TS \add_x_22_5/U132  ( .A(\add_x_22_5/n110 ), .B(\add_x_22_5/n109 ), 
        .Y(\add_x_22_5/n106 ) );
  NOR2X1TS \add_x_22_5/U127  ( .A(\add_x_22_5/n110 ), .B(\add_x_22_5/n103 ), 
        .Y(\add_x_22_5/n102 ) );
  NOR2X1TS \add_x_22_5/U21  ( .A(\add_x_22_5/n24 ), .B(\add_x_22_5/n17 ), .Y(
        \add_x_22_5/n16 ) );
  NOR2X1TS \add_x_22_5/U85  ( .A(\add_x_22_5/n76 ), .B(\add_x_22_5/n69 ), .Y(
        \add_x_22_5/n68 ) );
  NOR2X1TS \add_x_22_5/U63  ( .A(\add_x_22_5/n58 ), .B(\add_x_22_5/n51 ), .Y(
        \add_x_22_5/n50 ) );
  NOR2X1TS \add_x_22_5/U43  ( .A(\add_x_22_5/n42 ), .B(\add_x_22_5/n35 ), .Y(
        \add_x_22_5/n34 ) );
  NOR2X1TS \add_x_22_5/U6  ( .A(\add_x_22_5/n26 ), .B(\add_x_22_5/n5 ), .Y(
        \add_x_22_5/n4 ) );
  NOR2X1TS \add_x_22_5/U12  ( .A(\add_x_22_5/n17 ), .B(\add_x_22_5/n10 ), .Y(
        \add_x_22_5/n9 ) );
  NOR2X1TS \add_x_22_5/U54  ( .A(\add_x_22_5/n51 ), .B(\add_x_22_5/n44 ), .Y(
        \add_x_22_5/n43 ) );
  NOR2X1TS \add_x_22_5/U68  ( .A(\add_x_22_5/n58 ), .B(\add_x_22_5/n57 ), .Y(
        \add_x_22_5/n54 ) );
  NOR2X1TS \add_x_22_5/U138  ( .A(\add_x_22_5/n112 ), .B(\add_x_22_5/n119 ), 
        .Y(\add_x_22_5/n111 ) );
  NOR2X1TS \add_x_22_5/U96  ( .A(\add_x_22_5/n87 ), .B(\add_x_22_5/n78 ), .Y(
        \add_x_22_5/n77 ) );
  XNOR2X1TS \add_x_22_5/U146  ( .A(\add_x_22_5/n121 ), .B(n2578), .Y(
        \addr_calc/iir_write_calc/counter/N44 ) );
  XNOR2X1TS \add_x_22_5/U80  ( .A(\add_x_22_5/n68 ), .B(\add_x_22_5/n67 ), .Y(
        \addr_calc/iir_write_calc/counter/N57 ) );
  NAND2X1TS \add_x_22_5/U123  ( .A(\add_x_22_5/n102 ), .B(n2039), .Y(
        \add_x_22_5/n99 ) );
  XNOR2X1TS \add_x_22_5/U93  ( .A(\add_x_22_5/n81 ), .B(\add_x_22_5/n80 ), .Y(
        \addr_calc/iir_write_calc/counter/N54 ) );
  XNOR2X1TS \add_x_22_5/U126  ( .A(\add_x_22_5/n106 ), .B(n1937), .Y(
        \addr_calc/iir_write_calc/counter/N48 ) );
  XNOR2X1TS \add_x_22_5/U142  ( .A(\add_x_22_5/n118 ), .B(\add_x_22_5/n117 ), 
        .Y(\addr_calc/iir_write_calc/counter/N45 ) );
  NAND2X1TS \add_x_22_5/U90  ( .A(\add_x_22_5/n75 ), .B(n2044), .Y(
        \add_x_22_5/n72 ) );
  XNOR2X1TS \add_x_22_5/U122  ( .A(\add_x_22_5/n102 ), .B(\add_x_22_5/n101 ), 
        .Y(\addr_calc/iir_write_calc/counter/N49 ) );
  XNOR2X1TS \add_x_22_5/U111  ( .A(\add_x_22_5/n93 ), .B(\add_x_22_5/n92 ), 
        .Y(\addr_calc/iir_write_calc/counter/N51 ) );
  XNOR2X1TS \add_x_22_5/U89  ( .A(\add_x_22_5/n75 ), .B(\add_x_22_5/n74 ), .Y(
        \addr_calc/iir_write_calc/counter/N55 ) );
  XNOR2X1TS \add_x_22_5/U16  ( .A(\add_x_22_5/n16 ), .B(\add_x_22_5/n15 ), .Y(
        \addr_calc/iir_write_calc/counter/N69 ) );
  NAND2X1TS \add_x_22_5/U17  ( .A(\add_x_22_5/n16 ), .B(n2573), .Y(
        \add_x_22_5/n13 ) );
  NAND2X1TS \add_x_22_5/U26  ( .A(\add_x_22_5/n23 ), .B(
        \addr_calc/iir_write_calc/count[24] ), .Y(\add_x_22_5/n20 ) );
  XNOR2X1TS \add_x_22_5/U25  ( .A(\add_x_22_5/n23 ), .B(n2050), .Y(
        \addr_calc/iir_write_calc/counter/N67 ) );
  NAND2X1TS \add_x_22_5/U11  ( .A(\add_x_22_5/n23 ), .B(\add_x_22_5/n9 ), .Y(
        \add_x_22_5/n8 ) );
  NAND2X1TS \add_x_22_5/U39  ( .A(\add_x_22_5/n34 ), .B(n2579), .Y(
        \add_x_22_5/n31 ) );
  NAND2X1TS \add_x_22_5/U95  ( .A(\add_x_22_5/n93 ), .B(\add_x_22_5/n77 ), .Y(
        \add_x_22_5/n76 ) );
  NAND2X1TS \add_x_22_5/U59  ( .A(\add_x_22_5/n50 ), .B(n2571), .Y(
        \add_x_22_5/n47 ) );
  XNOR2X1TS \add_x_22_5/U38  ( .A(\add_x_22_5/n34 ), .B(\add_x_22_5/n33 ), .Y(
        \addr_calc/iir_write_calc/counter/N65 ) );
  NAND2X1TS \add_x_22_5/U53  ( .A(\add_x_22_5/n59 ), .B(\add_x_22_5/n43 ), .Y(
        \add_x_22_5/n42 ) );
  ADDHXLTS \add_x_22_5/U2  ( .A(n1854), .B(\add_x_22_5/n2 ), .CO(
        \add_x_22_5/n1 ), .S(\addr_calc/iir_write_calc/counter/N73 ) );
  NAND2X1TS \add_x_22_5/U5  ( .A(\add_x_22_5/n4 ), .B(\add_x_22_5/n59 ), .Y(
        \add_x_22_5/n3 ) );
  NAND2X1TS \add_x_22_5/U22  ( .A(n2051), .B(n1969), .Y(\add_x_22_5/n17 ) );
  NAND2X1TS \add_x_22_5/U44  ( .A(n2048), .B(n1962), .Y(\add_x_22_5/n35 ) );
  NAND2X1TS \add_x_22_5/U55  ( .A(n2571), .B(n1958), .Y(\add_x_22_5/n44 ) );
  NAND2X1TS \add_x_22_5/U64  ( .A(\addr_calc/iir_write_calc/count[16] ), .B(
        \addr_calc/iir_write_calc/count[17] ), .Y(\add_x_22_5/n51 ) );
  XNOR2X1TS \add_x_22_5/U62  ( .A(\add_x_22_5/n54 ), .B(\add_x_22_5/n53 ), .Y(
        \addr_calc/iir_write_calc/counter/N60 ) );
  NAND2X1TS \add_x_22_5/U148  ( .A(n1931), .B(
        \addr_calc/iir_write_calc/count[0] ), .Y(\add_x_22_5/n119 ) );
  NAND2X1TS \add_x_22_5/U139  ( .A(n2036), .B(n1933), .Y(\add_x_22_5/n112 ) );
  NAND2X1TS \add_x_22_5/U128  ( .A(\addr_calc/iir_write_calc/count[4] ), .B(
        \addr_calc/iir_write_calc/count[5] ), .Y(\add_x_22_5/n103 ) );
  NAND2X1TS \add_x_22_5/U86  ( .A(\addr_calc/iir_write_calc/count[12] ), .B(
        \addr_calc/iir_write_calc/count[13] ), .Y(\add_x_22_5/n69 ) );
  NAND2X1TS \add_x_22_5/U97  ( .A(\addr_calc/iir_write_calc/count[10] ), .B(
        \addr_calc/iir_write_calc/count[11] ), .Y(\add_x_22_5/n78 ) );
  NAND2X1TS \add_x_22_5/U108  ( .A(\addr_calc/iir_write_calc/count[8] ), .B(
        \addr_calc/iir_write_calc/count[9] ), .Y(\add_x_22_5/n87 ) );
  XOR2X1TS \add_x_22_5/U136  ( .A(\add_x_22_5/n115 ), .B(\add_x_22_5/n114 ), 
        .Y(\addr_calc/iir_write_calc/counter/N46 ) );
  XOR2X1TS \add_x_22_5/U131  ( .A(\add_x_22_5/n110 ), .B(\add_x_22_5/n109 ), 
        .Y(\addr_calc/iir_write_calc/counter/N47 ) );
  XOR2X1TS \add_x_22_5/U115  ( .A(\add_x_22_5/n99 ), .B(n1938), .Y(
        \addr_calc/iir_write_calc/counter/N50 ) );
  XOR2X1TS \add_x_22_5/U105  ( .A(\add_x_22_5/n90 ), .B(\add_x_22_5/n89 ), .Y(
        \addr_calc/iir_write_calc/counter/N52 ) );
  XOR2X1TS \add_x_22_5/U100  ( .A(\add_x_22_5/n85 ), .B(\add_x_22_5/n84 ), .Y(
        \addr_calc/iir_write_calc/counter/N53 ) );
  XOR2X1TS \add_x_22_5/U84  ( .A(\add_x_22_5/n72 ), .B(\add_x_22_5/n71 ), .Y(
        \addr_calc/iir_write_calc/counter/N56 ) );
  XOR2X1TS \add_x_22_5/U51  ( .A(\add_x_22_5/n47 ), .B(n1957), .Y(
        \addr_calc/iir_write_calc/counter/N62 ) );
  XOR2X1TS \add_x_22_5/U29  ( .A(\add_x_22_5/n31 ), .B(n1964), .Y(
        \addr_calc/iir_write_calc/counter/N66 ) );
  XOR2X1TS \add_x_22_5/U20  ( .A(\add_x_22_5/n20 ), .B(n1968), .Y(
        \addr_calc/iir_write_calc/counter/N68 ) );
  XOR2X1TS \add_x_22_5/U10  ( .A(\add_x_22_5/n13 ), .B(n1971), .Y(
        \addr_calc/iir_write_calc/counter/N70 ) );
  XOR2X1TS \add_x_22_5/U4  ( .A(\add_x_22_5/n8 ), .B(n1973), .Y(
        \addr_calc/iir_write_calc/counter/N71 ) );
  AHHCINX2TS \add_x_22_5/U3  ( .A(n1851), .CIN(\add_x_22_5/n3 ), .S(
        \addr_calc/iir_write_calc/counter/N72 ), .CO(\add_x_22_5/n2 ) );
  XOR2X1TS \add_x_22_5/U1  ( .A(\add_x_22_5/n1 ), .B(n1857), .Y(
        \addr_calc/iir_write_calc/counter/N74 ) );
  NOR2X1TS \add_x_22_3/U101  ( .A(\add_x_22_3/n85 ), .B(\add_x_22_3/n84 ), .Y(
        \add_x_22_3/n81 ) );
  NOR2X1TS \add_x_22_3/U132  ( .A(\add_x_22_3/n110 ), .B(\add_x_22_3/n109 ), 
        .Y(\add_x_22_3/n106 ) );
  NOR2X1TS \add_x_22_3/U127  ( .A(\add_x_22_3/n110 ), .B(\add_x_22_3/n103 ), 
        .Y(\add_x_22_3/n102 ) );
  NOR2X1TS \add_x_22_3/U63  ( .A(\add_x_22_3/n58 ), .B(\add_x_22_3/n51 ), .Y(
        \add_x_22_3/n50 ) );
  NOR2X1TS \add_x_22_3/U85  ( .A(\add_x_22_3/n76 ), .B(\add_x_22_3/n69 ), .Y(
        \add_x_22_3/n68 ) );
  NOR2X1TS \add_x_22_3/U43  ( .A(\add_x_22_3/n42 ), .B(\add_x_22_3/n35 ), .Y(
        \add_x_22_3/n34 ) );
  NOR2X1TS \add_x_22_3/U21  ( .A(\add_x_22_3/n24 ), .B(\add_x_22_3/n17 ), .Y(
        \add_x_22_3/n16 ) );
  NOR2X1TS \add_x_22_3/U12  ( .A(\add_x_22_3/n17 ), .B(\add_x_22_3/n10 ), .Y(
        \add_x_22_3/n9 ) );
  NOR2X1TS \add_x_22_3/U34  ( .A(\add_x_22_3/n35 ), .B(\add_x_22_3/n28 ), .Y(
        \add_x_22_3/n27 ) );
  NOR2X1TS \add_x_22_3/U54  ( .A(\add_x_22_3/n51 ), .B(\add_x_22_3/n44 ), .Y(
        \add_x_22_3/n43 ) );
  NOR2X1TS \add_x_22_3/U68  ( .A(\add_x_22_3/n58 ), .B(\add_x_22_3/n57 ), .Y(
        \add_x_22_3/n54 ) );
  NOR2X1TS \add_x_22_3/U138  ( .A(\add_x_22_3/n112 ), .B(\add_x_22_3/n119 ), 
        .Y(\add_x_22_3/n111 ) );
  NOR2X1TS \add_x_22_3/U96  ( .A(\add_x_22_3/n87 ), .B(\add_x_22_3/n78 ), .Y(
        \add_x_22_3/n77 ) );
  XNOR2X1TS \add_x_22_3/U142  ( .A(\add_x_22_3/n118 ), .B(n1989), .Y(
        \addr_calc/fir_write_calc/counter/N45 ) );
  NAND2X1TS \add_x_22_3/U143  ( .A(\add_x_22_3/n118 ), .B(
        \addr_calc/fir_write_calc/count[2] ), .Y(\add_x_22_3/n115 ) );
  XNOR2X1TS \add_x_22_3/U111  ( .A(\add_x_22_3/n93 ), .B(\add_x_22_3/n92 ), 
        .Y(\addr_calc/fir_write_calc/counter/N51 ) );
  XNOR2X1TS \add_x_22_3/U93  ( .A(\add_x_22_3/n81 ), .B(\add_x_22_3/n80 ), .Y(
        \addr_calc/fir_write_calc/counter/N54 ) );
  XNOR2X1TS \add_x_22_3/U126  ( .A(\add_x_22_3/n106 ), .B(\add_x_22_3/n105 ), 
        .Y(\addr_calc/fir_write_calc/counter/N48 ) );
  XNOR2X1TS \add_x_22_3/U38  ( .A(\add_x_22_3/n34 ), .B(n2012), .Y(
        \addr_calc/fir_write_calc/counter/N65 ) );
  XNOR2X1TS \add_x_22_3/U122  ( .A(\add_x_22_3/n102 ), .B(\add_x_22_3/n101 ), 
        .Y(\addr_calc/fir_write_calc/counter/N49 ) );
  XNOR2X1TS \add_x_22_3/U80  ( .A(\add_x_22_3/n68 ), .B(n2002), .Y(
        \addr_calc/fir_write_calc/counter/N57 ) );
  XNOR2X1TS \add_x_22_3/U58  ( .A(\add_x_22_3/n50 ), .B(n2005), .Y(
        \addr_calc/fir_write_calc/counter/N61 ) );
  NAND2X1TS \add_x_22_3/U90  ( .A(\add_x_22_3/n75 ), .B(n2000), .Y(
        \add_x_22_3/n72 ) );
  NAND2X1TS \add_x_22_3/U59  ( .A(\add_x_22_3/n50 ), .B(n2006), .Y(
        \add_x_22_3/n47 ) );
  NAND2X1TS \add_x_22_3/U95  ( .A(\add_x_22_3/n93 ), .B(\add_x_22_3/n77 ), .Y(
        \add_x_22_3/n76 ) );
  NAND2X1TS \add_x_22_3/U17  ( .A(\add_x_22_3/n16 ), .B(n2581), .Y(
        \add_x_22_3/n13 ) );
  NAND2X1TS \add_x_22_3/U39  ( .A(\add_x_22_3/n34 ), .B(n1668), .Y(
        \add_x_22_3/n31 ) );
  NAND2X1TS \add_x_22_3/U53  ( .A(\add_x_22_3/n59 ), .B(\add_x_22_3/n43 ), .Y(
        \add_x_22_3/n42 ) );
  NAND2X1TS \add_x_22_3/U11  ( .A(\add_x_22_3/n23 ), .B(\add_x_22_3/n9 ), .Y(
        \add_x_22_3/n8 ) );
  ADDHXLTS \add_x_22_3/U2  ( .A(n1836), .B(\add_x_22_3/n2 ), .CO(
        \add_x_22_3/n1 ), .S(\addr_calc/fir_write_calc/counter/N73 ) );
  NAND2X1TS \add_x_22_3/U22  ( .A(n2577), .B(n1894), .Y(\add_x_22_3/n17 ) );
  NAND2X1TS \add_x_22_3/U26  ( .A(\add_x_22_3/n23 ), .B(n2577), .Y(
        \add_x_22_3/n20 ) );
  XNOR2X1TS \add_x_22_3/U25  ( .A(\add_x_22_3/n23 ), .B(\add_x_22_3/n22 ), .Y(
        \addr_calc/fir_write_calc/counter/N67 ) );
  NAND2X1TS \add_x_22_3/U33  ( .A(\add_x_22_3/n43 ), .B(\add_x_22_3/n27 ), .Y(
        \add_x_22_3/n26 ) );
  NAND2X1TS \add_x_22_3/U44  ( .A(n1669), .B(n1892), .Y(\add_x_22_3/n35 ) );
  NAND2X1TS \add_x_22_3/U55  ( .A(n2006), .B(n1670), .Y(\add_x_22_3/n44 ) );
  NAND2X1TS \add_x_22_3/U64  ( .A(n2564), .B(
        \addr_calc/fir_write_calc/count[17] ), .Y(\add_x_22_3/n51 ) );
  XNOR2X1TS \add_x_22_3/U62  ( .A(\add_x_22_3/n54 ), .B(n1885), .Y(
        \addr_calc/fir_write_calc/counter/N60 ) );
  NAND2X1TS \add_x_22_3/U148  ( .A(\addr_calc/fir_write_calc/count[1] ), .B(
        \addr_calc/fir_write_calc/count[0] ), .Y(\add_x_22_3/n119 ) );
  NAND2X1TS \add_x_22_3/U139  ( .A(n1990), .B(
        \addr_calc/fir_write_calc/count[3] ), .Y(\add_x_22_3/n112 ) );
  NAND2X1TS \add_x_22_3/U128  ( .A(\addr_calc/fir_write_calc/count[4] ), .B(
        n1867), .Y(\add_x_22_3/n103 ) );
  NAND2X1TS \add_x_22_3/U86  ( .A(n1999), .B(n1880), .Y(\add_x_22_3/n69 ) );
  NAND2X1TS \add_x_22_3/U97  ( .A(n1874), .B(
        \addr_calc/fir_write_calc/count[11] ), .Y(\add_x_22_3/n78 ) );
  NAND2X1TS \add_x_22_3/U108  ( .A(n1995), .B(
        \addr_calc/fir_write_calc/count[9] ), .Y(\add_x_22_3/n87 ) );
  XOR2X1TS \add_x_22_3/U136  ( .A(\add_x_22_3/n115 ), .B(\add_x_22_3/n114 ), 
        .Y(\addr_calc/fir_write_calc/counter/N46 ) );
  XOR2X1TS \add_x_22_3/U105  ( .A(\add_x_22_3/n90 ), .B(\add_x_22_3/n89 ), .Y(
        \addr_calc/fir_write_calc/counter/N52 ) );
  XOR2X1TS \add_x_22_3/U84  ( .A(\add_x_22_3/n72 ), .B(\add_x_22_3/n71 ), .Y(
        \addr_calc/fir_write_calc/counter/N56 ) );
  XOR2X1TS \add_x_22_3/U67  ( .A(\add_x_22_3/n58 ), .B(\add_x_22_3/n57 ), .Y(
        \addr_calc/fir_write_calc/counter/N59 ) );
  XOR2X1TS \add_x_22_3/U51  ( .A(\add_x_22_3/n47 ), .B(n1889), .Y(
        \addr_calc/fir_write_calc/counter/N62 ) );
  XOR2X1TS \add_x_22_3/U29  ( .A(\add_x_22_3/n31 ), .B(\add_x_22_3/n30 ), .Y(
        \addr_calc/fir_write_calc/counter/N66 ) );
  XOR2X1TS \add_x_22_3/U20  ( .A(\add_x_22_3/n20 ), .B(\add_x_22_3/n19 ), .Y(
        \addr_calc/fir_write_calc/counter/N68 ) );
  XOR2X1TS \add_x_22_3/U10  ( .A(\add_x_22_3/n13 ), .B(n1834), .Y(
        \addr_calc/fir_write_calc/counter/N70 ) );
  XOR2X1TS \add_x_22_3/U4  ( .A(\add_x_22_3/n8 ), .B(\add_x_22_3/n7 ), .Y(
        \addr_calc/fir_write_calc/counter/N71 ) );
  XOR2X1TS \add_x_22_3/U1  ( .A(\add_x_22_3/n1 ), .B(n2550), .Y(
        \addr_calc/fir_write_calc/counter/N74 ) );
  NOR2X1TS \add_x_22_2/U68  ( .A(\add_x_22_2/n58 ), .B(n1887), .Y(
        \add_x_22_2/n54 ) );
  NOR2X1TS \add_x_22_2/U127  ( .A(\add_x_22_2/n110 ), .B(\add_x_22_2/n103 ), 
        .Y(\add_x_22_2/n102 ) );
  NOR2X1TS \add_x_22_2/U101  ( .A(\add_x_22_2/n85 ), .B(n1897), .Y(
        \add_x_22_2/n81 ) );
  NOR2X1TS \add_x_22_2/U85  ( .A(\add_x_22_2/n76 ), .B(\add_x_22_2/n69 ), .Y(
        \add_x_22_2/n68 ) );
  NOR2X1TS \add_x_22_2/U63  ( .A(\add_x_22_2/n58 ), .B(\add_x_22_2/n51 ), .Y(
        \add_x_22_2/n50 ) );
  NOR2X1TS \add_x_22_2/U43  ( .A(\add_x_22_2/n42 ), .B(\add_x_22_2/n35 ), .Y(
        \add_x_22_2/n34 ) );
  NOR2X1TS \add_x_22_2/U12  ( .A(\add_x_22_2/n17 ), .B(\add_x_22_2/n10 ), .Y(
        \add_x_22_2/n9 ) );
  NOR2X1TS \add_x_22_2/U21  ( .A(\add_x_22_2/n24 ), .B(\add_x_22_2/n17 ), .Y(
        \add_x_22_2/n16 ) );
  NOR2X1TS \add_x_22_2/U54  ( .A(\add_x_22_2/n51 ), .B(\add_x_22_2/n44 ), .Y(
        \add_x_22_2/n43 ) );
  NOR2X1TS \add_x_22_2/U138  ( .A(\add_x_22_2/n112 ), .B(\add_x_22_2/n119 ), 
        .Y(\add_x_22_2/n111 ) );
  NOR2X1TS \add_x_22_2/U96  ( .A(\add_x_22_2/n87 ), .B(\add_x_22_2/n78 ), .Y(
        \add_x_22_2/n77 ) );
  XNOR2X1TS \add_x_22_2/U142  ( .A(\add_x_22_2/n118 ), .B(\add_x_22_2/n117 ), 
        .Y(\addr_calc/fir_read_calc/counter/N45 ) );
  XNOR2X1TS \add_x_22_2/U58  ( .A(\add_x_22_2/n50 ), .B(n1987), .Y(
        \addr_calc/fir_read_calc/counter/N61 ) );
  XNOR2X1TS \add_x_22_2/U89  ( .A(\add_x_22_2/n75 ), .B(\add_x_22_2/n74 ), .Y(
        \addr_calc/fir_read_calc/counter/N55 ) );
  XNOR2X1TS \add_x_22_2/U122  ( .A(\add_x_22_2/n102 ), .B(\add_x_22_2/n101 ), 
        .Y(\addr_calc/fir_read_calc/counter/N49 ) );
  XNOR2X1TS \add_x_22_2/U62  ( .A(\add_x_22_2/n54 ), .B(\add_x_22_2/n53 ), .Y(
        \addr_calc/fir_read_calc/counter/N60 ) );
  XNOR2X1TS \add_x_22_2/U126  ( .A(\add_x_22_2/n106 ), .B(\add_x_22_2/n105 ), 
        .Y(\addr_calc/fir_read_calc/counter/N48 ) );
  XNOR2X1TS \add_x_22_2/U47  ( .A(\add_x_22_2/n41 ), .B(n1984), .Y(
        \addr_calc/fir_read_calc/counter/N63 ) );
  NAND2X1TS \add_x_22_2/U90  ( .A(\add_x_22_2/n75 ), .B(n1994), .Y(
        \add_x_22_2/n72 ) );
  XNOR2X1TS \add_x_22_2/U80  ( .A(\add_x_22_2/n68 ), .B(n1991), .Y(
        \addr_calc/fir_read_calc/counter/N57 ) );
  NAND2X1TS \add_x_22_2/U48  ( .A(\add_x_22_2/n41 ), .B(
        \addr_calc/fir_read_calc/count[20] ), .Y(\add_x_22_2/n38 ) );
  XNOR2X1TS \add_x_22_2/U93  ( .A(\add_x_22_2/n81 ), .B(\add_x_22_2/n80 ), .Y(
        \addr_calc/fir_read_calc/counter/N54 ) );
  NAND2X1TS \add_x_22_2/U95  ( .A(\add_x_22_2/n93 ), .B(\add_x_22_2/n77 ), .Y(
        \add_x_22_2/n76 ) );
  XNOR2X1TS \add_x_22_2/U38  ( .A(\add_x_22_2/n34 ), .B(n1981), .Y(
        \addr_calc/fir_read_calc/counter/N65 ) );
  XNOR2X1TS \add_x_22_2/U111  ( .A(\add_x_22_2/n93 ), .B(\add_x_22_2/n92 ), 
        .Y(\addr_calc/fir_read_calc/counter/N51 ) );
  NAND2X1TS \add_x_22_2/U59  ( .A(\add_x_22_2/n50 ), .B(
        \addr_calc/fir_read_calc/count[18] ), .Y(\add_x_22_2/n47 ) );
  XNOR2X1TS \add_x_22_2/U25  ( .A(\add_x_22_2/n23 ), .B(n1982), .Y(
        \addr_calc/fir_read_calc/counter/N67 ) );
  NAND2X1TS \add_x_22_2/U39  ( .A(\add_x_22_2/n34 ), .B(n1691), .Y(
        \add_x_22_2/n31 ) );
  NAND2X1TS \add_x_22_2/U53  ( .A(\add_x_22_2/n59 ), .B(\add_x_22_2/n43 ), .Y(
        \add_x_22_2/n42 ) );
  ADDHXLTS \add_x_22_2/U2  ( .A(\addr_calc/fir_read_calc/count[30] ), .B(
        \add_x_22_2/n2 ), .CO(\add_x_22_2/n1 ), .S(
        \addr_calc/fir_read_calc/counter/N73 ) );
  NAND2X1TS \add_x_22_2/U11  ( .A(\add_x_22_2/n23 ), .B(\add_x_22_2/n9 ), .Y(
        \add_x_22_2/n8 ) );
  NAND2X1TS \add_x_22_2/U22  ( .A(\addr_calc/fir_read_calc/count[24] ), .B(
        \addr_calc/fir_read_calc/count[25] ), .Y(\add_x_22_2/n17 ) );
  NAND2X1TS \add_x_22_2/U44  ( .A(\addr_calc/fir_read_calc/count[20] ), .B(
        n1879), .Y(\add_x_22_2/n35 ) );
  NAND2X1TS \add_x_22_2/U55  ( .A(\addr_calc/fir_read_calc/count[18] ), .B(
        n1881), .Y(\add_x_22_2/n44 ) );
  NAND2X1TS \add_x_22_2/U64  ( .A(n1888), .B(n1884), .Y(\add_x_22_2/n51 ) );
  NAND2X1TS \add_x_22_2/U148  ( .A(\addr_calc/fir_read_calc/count[1] ), .B(
        \addr_calc/fir_read_calc/count[0] ), .Y(\add_x_22_2/n119 ) );
  NAND2X1TS \add_x_22_2/U139  ( .A(\addr_calc/fir_read_calc/count[2] ), .B(
        \addr_calc/fir_read_calc/count[3] ), .Y(\add_x_22_2/n112 ) );
  NAND2X1TS \add_x_22_2/U128  ( .A(n1906), .B(
        \addr_calc/fir_read_calc/count[5] ), .Y(\add_x_22_2/n103 ) );
  NAND2X1TS \add_x_22_2/U86  ( .A(\addr_calc/fir_read_calc/count[12] ), .B(
        n1893), .Y(\add_x_22_2/n69 ) );
  NAND2X1TS \add_x_22_2/U97  ( .A(n1540), .B(
        \addr_calc/fir_read_calc/count[11] ), .Y(\add_x_22_2/n78 ) );
  NAND2X1TS \add_x_22_2/U108  ( .A(\addr_calc/fir_read_calc/count[8] ), .B(
        n1900), .Y(\add_x_22_2/n87 ) );
  XOR2X1TS \add_x_22_2/U131  ( .A(\add_x_22_2/n110 ), .B(\add_x_22_2/n109 ), 
        .Y(\addr_calc/fir_read_calc/counter/N47 ) );
  XOR2X1TS \add_x_22_2/U115  ( .A(\add_x_22_2/n99 ), .B(\add_x_22_2/n98 ), .Y(
        \addr_calc/fir_read_calc/counter/N50 ) );
  XOR2X1TS \add_x_22_2/U105  ( .A(\add_x_22_2/n90 ), .B(n1899), .Y(
        \addr_calc/fir_read_calc/counter/N52 ) );
  XOR2X1TS \add_x_22_2/U100  ( .A(\add_x_22_2/n85 ), .B(n1897), .Y(
        \addr_calc/fir_read_calc/counter/N53 ) );
  XOR2X1TS \add_x_22_2/U84  ( .A(\add_x_22_2/n72 ), .B(\add_x_22_2/n71 ), .Y(
        \addr_calc/fir_read_calc/counter/N56 ) );
  XOR2X1TS \add_x_22_2/U67  ( .A(\add_x_22_2/n58 ), .B(n1887), .Y(
        \addr_calc/fir_read_calc/counter/N59 ) );
  XOR2X1TS \add_x_22_2/U51  ( .A(\add_x_22_2/n47 ), .B(\add_x_22_2/n46 ), .Y(
        \addr_calc/fir_read_calc/counter/N62 ) );
  XOR2X1TS \add_x_22_2/U42  ( .A(\add_x_22_2/n38 ), .B(n1878), .Y(
        \addr_calc/fir_read_calc/counter/N64 ) );
  XOR2X1TS \add_x_22_2/U29  ( .A(\add_x_22_2/n31 ), .B(\add_x_22_2/n30 ), .Y(
        \addr_calc/fir_read_calc/counter/N66 ) );
  XOR2X1TS \add_x_22_2/U4  ( .A(\add_x_22_2/n8 ), .B(n1870), .Y(
        \addr_calc/fir_read_calc/counter/N71 ) );
  NOR2X1TS \add_x_22_0/U127  ( .A(\add_x_22_0/n110 ), .B(\add_x_22_0/n103 ), 
        .Y(\add_x_22_0/n102 ) );
  NOR2X1TS \add_x_22_0/U132  ( .A(\add_x_22_0/n110 ), .B(\add_x_22_0/n109 ), 
        .Y(\add_x_22_0/n106 ) );
  NOR2X1TS \add_x_22_0/U85  ( .A(\add_x_22_0/n76 ), .B(\add_x_22_0/n69 ), .Y(
        \add_x_22_0/n68 ) );
  NOR2X1TS \add_x_22_0/U21  ( .A(\add_x_22_0/n24 ), .B(\add_x_22_0/n17 ), .Y(
        \add_x_22_0/n16 ) );
  NOR2X1TS \add_x_22_0/U43  ( .A(\add_x_22_0/n42 ), .B(\add_x_22_0/n35 ), .Y(
        \add_x_22_0/n34 ) );
  NOR2X1TS \add_x_22_0/U6  ( .A(\add_x_22_0/n26 ), .B(\add_x_22_0/n5 ), .Y(
        \add_x_22_0/n4 ) );
  NOR2X1TS \add_x_22_0/U12  ( .A(\add_x_22_0/n17 ), .B(\add_x_22_0/n10 ), .Y(
        \add_x_22_0/n9 ) );
  NOR2X1TS \add_x_22_0/U54  ( .A(\add_x_22_0/n51 ), .B(\add_x_22_0/n44 ), .Y(
        \add_x_22_0/n43 ) );
  NOR2X1TS \add_x_22_0/U63  ( .A(\add_x_22_0/n58 ), .B(\add_x_22_0/n51 ), .Y(
        \add_x_22_0/n50 ) );
  NOR2X1TS \add_x_22_0/U138  ( .A(\add_x_22_0/n112 ), .B(\add_x_22_0/n119 ), 
        .Y(\add_x_22_0/n111 ) );
  NOR2X1TS \add_x_22_0/U118  ( .A(\add_x_22_0/n103 ), .B(\add_x_22_0/n96 ), 
        .Y(\add_x_22_0/n95 ) );
  NOR2X1TS \add_x_22_0/U96  ( .A(\add_x_22_0/n87 ), .B(\add_x_22_0/n78 ), .Y(
        \add_x_22_0/n77 ) );
  XNOR2X1TS \add_x_22_0/U146  ( .A(\add_x_22_0/n121 ), .B(
        \addr_calc/fft_read_calc/count[0] ), .Y(
        \addr_calc/fft_read_calc/counter/N44 ) );
  XNOR2X1TS \add_x_22_0/U142  ( .A(\add_x_22_0/n118 ), .B(\add_x_22_0/n117 ), 
        .Y(\addr_calc/fft_read_calc/counter/N45 ) );
  XNOR2X1TS \add_x_22_0/U89  ( .A(\add_x_22_0/n75 ), .B(n2045), .Y(
        \addr_calc/fft_read_calc/counter/N55 ) );
  XNOR2X1TS \add_x_22_0/U47  ( .A(\add_x_22_0/n41 ), .B(\add_x_22_0/n40 ), .Y(
        \addr_calc/fft_read_calc/counter/N63 ) );
  NAND2X1TS \add_x_22_0/U143  ( .A(\add_x_22_0/n118 ), .B(n2056), .Y(
        \add_x_22_0/n115 ) );
  XNOR2X1TS \add_x_22_0/U80  ( .A(\add_x_22_0/n68 ), .B(n2042), .Y(
        \addr_calc/fft_read_calc/counter/N57 ) );
  XNOR2X1TS \add_x_22_0/U38  ( .A(\add_x_22_0/n34 ), .B(n2040), .Y(
        \addr_calc/fft_read_calc/counter/N65 ) );
  XNOR2X1TS \add_x_22_0/U111  ( .A(\add_x_22_0/n93 ), .B(\add_x_22_0/n92 ), 
        .Y(\addr_calc/fft_read_calc/counter/N51 ) );
  NAND2X1TS \add_x_22_0/U90  ( .A(\add_x_22_0/n75 ), .B(
        \addr_calc/fft_read_calc/count[12] ), .Y(\add_x_22_0/n72 ) );
  XNOR2X1TS \add_x_22_0/U126  ( .A(\add_x_22_0/n106 ), .B(\add_x_22_0/n105 ), 
        .Y(\addr_calc/fft_read_calc/counter/N48 ) );
  NAND2X1TS \add_x_22_0/U95  ( .A(\add_x_22_0/n93 ), .B(\add_x_22_0/n77 ), .Y(
        \add_x_22_0/n76 ) );
  NAND2X1TS \add_x_22_0/U26  ( .A(\add_x_22_0/n23 ), .B(
        \addr_calc/fft_read_calc/count[24] ), .Y(\add_x_22_0/n20 ) );
  NAND2X1TS \add_x_22_0/U11  ( .A(\add_x_22_0/n23 ), .B(\add_x_22_0/n9 ), .Y(
        \add_x_22_0/n8 ) );
  NAND2X1TS \add_x_22_0/U17  ( .A(\add_x_22_0/n16 ), .B(n2575), .Y(
        \add_x_22_0/n13 ) );
  NAND2X1TS \add_x_22_0/U39  ( .A(\add_x_22_0/n34 ), .B(n1665), .Y(
        \add_x_22_0/n31 ) );
  NAND2X1TS \add_x_22_0/U53  ( .A(\add_x_22_0/n59 ), .B(\add_x_22_0/n43 ), .Y(
        \add_x_22_0/n42 ) );
  XNOR2X1TS \add_x_22_0/U25  ( .A(\add_x_22_0/n23 ), .B(n2037), .Y(
        \addr_calc/fft_read_calc/counter/N67 ) );
  ADDHXLTS \add_x_22_0/U2  ( .A(\addr_calc/fft_read_calc/count[30] ), .B(
        \add_x_22_0/n2 ), .CO(\add_x_22_0/n1 ), .S(
        \addr_calc/fft_read_calc/counter/N73 ) );
  NAND2X1TS \add_x_22_0/U5  ( .A(\add_x_22_0/n4 ), .B(\add_x_22_0/n59 ), .Y(
        \add_x_22_0/n3 ) );
  NAND2X1TS \add_x_22_0/U7  ( .A(\add_x_22_0/n9 ), .B(n2559), .Y(
        \add_x_22_0/n5 ) );
  NAND2X1TS \add_x_22_0/U22  ( .A(\addr_calc/fft_read_calc/count[24] ), .B(
        \addr_calc/fft_read_calc/count[25] ), .Y(\add_x_22_0/n17 ) );
  NAND2X1TS \add_x_22_0/U44  ( .A(n2572), .B(n1953), .Y(\add_x_22_0/n35 ) );
  NAND2X1TS \add_x_22_0/U55  ( .A(n2569), .B(
        \addr_calc/fft_read_calc/count[19] ), .Y(\add_x_22_0/n44 ) );
  NAND2X1TS \add_x_22_0/U59  ( .A(\add_x_22_0/n50 ), .B(n2569), .Y(
        \add_x_22_0/n47 ) );
  NAND2X1TS \add_x_22_0/U64  ( .A(n2554), .B(
        \addr_calc/fft_read_calc/count[17] ), .Y(\add_x_22_0/n51 ) );
  NAND2X1TS \add_x_22_0/U117  ( .A(\add_x_22_0/n95 ), .B(\add_x_22_0/n111 ), 
        .Y(\add_x_22_0/n94 ) );
  NAND2X1TS \add_x_22_0/U148  ( .A(n1979), .B(n2058), .Y(\add_x_22_0/n119 ) );
  NAND2X1TS \add_x_22_0/U139  ( .A(n2056), .B(
        \addr_calc/fft_read_calc/count[3] ), .Y(\add_x_22_0/n112 ) );
  NAND2X1TS \add_x_22_0/U119  ( .A(n2052), .B(
        \addr_calc/fft_read_calc/count[7] ), .Y(\add_x_22_0/n96 ) );
  NAND2X1TS \add_x_22_0/U128  ( .A(n2552), .B(n1977), .Y(\add_x_22_0/n103 ) );
  NAND2X1TS \add_x_22_0/U86  ( .A(n2046), .B(n1967), .Y(\add_x_22_0/n69 ) );
  NAND2X1TS \add_x_22_0/U97  ( .A(\addr_calc/fft_read_calc/count[10] ), .B(
        \addr_calc/fft_read_calc/count[11] ), .Y(\add_x_22_0/n78 ) );
  NAND2X1TS \add_x_22_0/U108  ( .A(\addr_calc/fft_read_calc/count[8] ), .B(
        \addr_calc/fft_read_calc/count[9] ), .Y(\add_x_22_0/n87 ) );
  XOR2X1TS \add_x_22_0/U136  ( .A(\add_x_22_0/n115 ), .B(\add_x_22_0/n114 ), 
        .Y(\addr_calc/fft_read_calc/counter/N46 ) );
  XOR2X1TS \add_x_22_0/U115  ( .A(\add_x_22_0/n99 ), .B(n1975), .Y(
        \addr_calc/fft_read_calc/counter/N50 ) );
  XOR2X1TS \add_x_22_0/U105  ( .A(\add_x_22_0/n90 ), .B(\add_x_22_0/n89 ), .Y(
        \addr_calc/fft_read_calc/counter/N52 ) );
  XOR2X1TS \add_x_22_0/U100  ( .A(\add_x_22_0/n85 ), .B(\add_x_22_0/n84 ), .Y(
        \addr_calc/fft_read_calc/counter/N53 ) );
  XOR2X1TS \add_x_22_0/U84  ( .A(\add_x_22_0/n72 ), .B(n1966), .Y(
        \addr_calc/fft_read_calc/counter/N56 ) );
  XOR2X1TS \add_x_22_0/U72  ( .A(\add_x_22_0/n65 ), .B(n1963), .Y(
        \addr_calc/fft_read_calc/counter/N58 ) );
  XOR2X1TS \add_x_22_0/U51  ( .A(\add_x_22_0/n47 ), .B(n1955), .Y(
        \addr_calc/fft_read_calc/counter/N62 ) );
  XOR2X1TS \add_x_22_0/U29  ( .A(\add_x_22_0/n31 ), .B(n1949), .Y(
        \addr_calc/fft_read_calc/counter/N66 ) );
  XOR2X1TS \add_x_22_0/U20  ( .A(\add_x_22_0/n20 ), .B(n1946), .Y(
        \addr_calc/fft_read_calc/counter/N68 ) );
  XOR2X1TS \add_x_22_0/U10  ( .A(\add_x_22_0/n13 ), .B(n1943), .Y(
        \addr_calc/fft_read_calc/counter/N70 ) );
  XOR2X1TS \add_x_22_0/U4  ( .A(\add_x_22_0/n8 ), .B(\add_x_22_0/n7 ), .Y(
        \addr_calc/fft_read_calc/counter/N71 ) );
  AHHCINX2TS \add_x_22_0/U3  ( .A(\addr_calc/fft_read_calc/count[29] ), .CIN(
        \add_x_22_0/n3 ), .S(\addr_calc/fft_read_calc/counter/N72 ), .CO(
        \add_x_22_0/n2 ) );
  DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[8]  ( .D(n963), .CK(clk), .Q(\addr_calc/iir_read_calc/count[8] ) );
  DFFHQX1TS \addr_calc/fir_read_calc/counter/count_reg[26]  ( .D(n1072), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[26] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[26]  ( .D(n1104), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[26] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[22]  ( .D(n980), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[22] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[24]  ( .D(n1106), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[24] ) );
  DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[26]  ( .D(n945), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[26] ) );
  DFFHQX1TS \addr_calc/fft_read_calc/counter/count_reg[26]  ( .D(n1008), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[26] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[26]  ( .D(n1040), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[26] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[26]  ( .D(n976), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[26] ) );
  DFFHQX1TS \addr_calc/iir_write_calc/counter/count_reg[18]  ( .D(n984), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[18] ) );
  DFFHQX1TS \addr_calc/iir_write_calc/counter/count_reg[14]  ( .D(n988), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[14] ) );
  DFFHQX1TS \addr_calc/fft_read_calc/counter/count_reg[18]  ( .D(n1016), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[18] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[3]  ( .D(n1063), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[3] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[16]  ( .D(n1050), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[16] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[16]  ( .D(n1114), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[16] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[23]  ( .D(n1107), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[23] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[9]  ( .D(n993), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[9] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[9]  ( .D(n1025), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[9] ) );
  DFFHQX1TS \addr_calc/fir_read_calc/counter/count_reg[23]  ( .D(n1075), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[23] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[28]  ( .D(n1038), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[28] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[23]  ( .D(n1043), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[23] ) );
  DFFHQX1TS \addr_calc/fft_read_calc/counter/count_reg[16]  ( .D(n1018), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[16] ) );
  DFFHQX1TS \addr_calc/fft_read_calc/counter/count_reg[4]  ( .D(n1030), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[4] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[31]  ( .D(n1099), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[31] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[31]  ( .D(n1132), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[31] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[2]  ( .D(n1032), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[2] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[8]  ( .D(n1026), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[8] ) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[12]  ( .D(n990), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[12] ) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[8]  ( .D(n994), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[8] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[0]  ( .D(n1066), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[0] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[2]  ( .D(n1064), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[2] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[8]  ( .D(n1058), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[8] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[12]  ( .D(n1054), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[12] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[14]  ( .D(n1052), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[14] ) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[6]  ( .D(n965), .CK(clk), .Q(\addr_calc/iir_read_calc/count[6] ) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[2]  ( .D(n969), .CK(clk), .Q(\addr_calc/iir_read_calc/count[2] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[2]  ( .D(n1096), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[2] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[6]  ( .D(n1092), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[6] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[8]  ( .D(n1090), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[8] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[8]  ( .D(n1122), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[8] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[12]  ( .D(n1086), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[12] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[6]  ( .D(n1124), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[6] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[0]  ( .D(n1130), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[0] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[1]  ( .D(n1033), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[1] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[3]  ( .D(n1031), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[3] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[5]  ( .D(n1029), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[5] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[10]  ( .D(n1024), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[10] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[11]  ( .D(n1023), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[11] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[1]  ( .D(n1065), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[1] ) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[10]  ( .D(n992), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[10] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[7]  ( .D(n1059), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[7] ) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[4]  ( .D(n998), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[4] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[9]  ( .D(n1057), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[9] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[3]  ( .D(n999), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[3] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[10]  ( .D(n1056), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[10] ) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[1]  ( .D(n1001), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[1] ) );
  DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[17]  ( .D(n1049), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[17] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[1]  ( .D(n1097), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[1] ) );
  DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[10]  ( .D(n961), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[10] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[3]  ( .D(n1095), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[3] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[4]  ( .D(n1094), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[4] ) );
  DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[7]  ( .D(n964), .CK(clk), .Q(\addr_calc/iir_read_calc/count[7] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[5]  ( .D(n1093), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[5] ) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[4]  ( .D(n967), .CK(clk), .Q(\addr_calc/iir_read_calc/count[4] ) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[1]  ( .D(n970), .CK(clk), .Q(\addr_calc/iir_read_calc/count[1] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[28]  ( .D(n1102), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[28] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[11]  ( .D(n1087), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[11] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[13]  ( .D(n1085), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[13] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[15]  ( .D(n1083), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[15] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[17]  ( .D(n1081), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[17] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[19]  ( .D(n1079), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[19] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[13]  ( .D(n1117), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[13] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[11]  ( .D(n1119), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[11] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[10]  ( .D(n1120), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[10] ) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[27]  ( .D(n1071), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[27] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[7]  ( .D(n1123), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[7] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[1]  ( .D(n1129), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[1] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[3]  ( .D(n1127), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[3] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[4]  ( .D(n1126), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[4] ) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[31]  ( .D(n1136), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[31] ) );
  DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[30]  ( .D(n1003), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[30] ) );
  DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[30]  ( .D(n1100), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[30] ) );
  TBUFX4TS \addr_calc/addr_tri6[13]  ( .A(\addr_calc/iir_write_addr[13] ), 
        .OE(n2779), .Y(addr[13]) );
  DFFQX2TS \addr_calc/iir_read_calc/counter/count_reg[12]  ( .D(n959), .CK(clk), .Q(\addr_calc/iir_read_calc/count[12] ) );
  DFFTRX2TS \addr_calc/fft_read_calc/counter/done_reg  ( .D(n783), .RN(n2072), 
        .CK(clk), .Q(fft_read_done), .QN(n895) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[28]  ( .D(n943), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[28] ) );
  DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[11]  ( .D(n960), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[11] ) );
  DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[13]  ( .D(n958), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[13] ) );
  TBUFX6TS \addr_calc/addr_tri5[18]  ( .A(\addr_calc/iir_read_addr[18] ), .OE(
        n2770), .Y(addr[18]) );
  DFFTRX2TS \addr_calc/iir_write_calc/counter/done_reg  ( .D(n787), .RN(
        iir_enable), .CK(clk), .Q(iir_write_done) );
  DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[19]  ( .D(n952), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[19] ) );
  DFFTRX2TS \addr_calc/fir_read_calc/counter/done_reg  ( .D(n1461), .RN(n2069), 
        .CK(clk), .Q(fir_read_done), .QN(n900) );
  DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[27]  ( .D(n944), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[27] ) );
  DFFQX2TS \addr_calc/iir_read_calc/counter/count_reg[31]  ( .D(n972), .CK(clk), .Q(\addr_calc/iir_read_calc/count[31] ) );
  DFFQX4TS \addr_calc/fft_read_calc/counter/count_reg[28]  ( .D(n1006), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[28] ) );
  DFFQX4TS \addr_calc/fft_read_calc/counter/count_reg[20]  ( .D(n1014), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[20] ) );
  DFFTRX2TS \addr_calc/fir_write_calc/counter/done_reg  ( .D(n785), .RN(
        fir_enable), .CK(clk), .Q(fir_write_done) );
  DFFHQX1TS \addr_calc/fir_write_calc/counter/count_reg[12]  ( .D(n1118), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[12] ) );
  DFFQX4TS \addr_calc/fir_write_calc/counter/count_reg[25]  ( .D(n1105), .CK(
        clk), .Q(\addr_calc/fir_write_calc/count[25] ) );
  AOI22XLTS U361 ( .A0(n2340), .A1(n2323), .B0(n2338), .B1(n2327), .Y(n930) );
  NAND2BXLTS U374 ( .AN(n2319), .B(n2334), .Y(n938) );
  NAND2XLTS \add_x_19_3/U5  ( .A(n2550), .B(n2381), .Y(\add_x_19_3/n34 ) );
  NAND2XLTS \DP_OP_158_296_6262/U1804  ( .A(\DP_OP_158_296_6262/n1837 ), .B(
        \DP_OP_158_296_6262/n1830 ), .Y(\DP_OP_158_296_6262/n1829 ) );
  NAND2XLTS \add_x_22_5/U13  ( .A(n2573), .B(
        \addr_calc/iir_write_calc/count[27] ), .Y(\add_x_22_5/n10 ) );
  NAND2XLTS \add_x_22_0/U13  ( .A(n2575), .B(
        \addr_calc/fft_read_calc/count[27] ), .Y(\add_x_22_0/n10 ) );
  NAND2XLTS \add_x_22_1/U13  ( .A(n2574), .B(
        \addr_calc/fft_write_calc/count[27] ), .Y(\add_x_22_1/n10 ) );
  NAND2XLTS \add_x_22_3/U13  ( .A(n2581), .B(
        \addr_calc/fir_write_calc/count[27] ), .Y(\add_x_22_3/n10 ) );
  NAND2XLTS \add_x_22_2/U13  ( .A(n2582), .B(n1873), .Y(\add_x_22_2/n10 ) );
  NOR2X1TS \add_x_19_0/U104  ( .A(n1956), .B(n2489), .Y(\add_x_19_0/n97 ) );
  OAI32X1TS U354 ( .A0(fir_read_done), .A1(n2071), .A2(fir_write_done), .B0(
        n2066), .B1(n2073), .Y(n928) );
  NAND2XLTS \add_x_19_0/U5  ( .A(\addr_calc/fft_read_calc/count[31] ), .B(
        n2382), .Y(\add_x_19_0/n34 ) );
  OAI21X1TS \add_x_19_5/U239  ( .A0(\add_x_19_5/n186 ), .A1(\add_x_19_5/n184 ), 
        .B0(\add_x_19_5/n185 ), .Y(\add_x_19_5/n183 ) );
  NOR3X1TS U356 ( .A(n1478), .B(fft_read_done), .C(n2587), .Y(n797) );
  NAND2X1TS \add_x_19_2/U67  ( .A(\add_x_19_2/n84 ), .B(\add_x_19_2/n76 ), .Y(
        \add_x_19_2/n74 ) );
  NAND2XLTS \add_x_22_5/U7  ( .A(\add_x_22_5/n9 ), .B(n1974), .Y(
        \add_x_22_5/n5 ) );
  NAND3XLTS U367 ( .A(n2069), .B(n934), .C(n2585), .Y(\data_cntl/N255 ) );
  AND2X2TS U389 ( .A(n2067), .B(n2585), .Y(n936) );
  NOR2X1TS \add_x_19_0/U24  ( .A(\add_x_19_0/n51 ), .B(\add_x_19_0/n48 ), .Y(
        \add_x_19_0/n46 ) );
  OAI211X1TS U348 ( .A0(n1829), .A1(n2059), .B0(iir_enable), .C0(n898), .Y(
        n926) );
  CLKINVX1TS U344 ( .A(n792), .Y(n923) );
  AOI211XLTS U363 ( .A0(n2340), .A1(n931), .B0(n2338), .C0(n932), .Y(
        \data_cntl/N257 ) );
  NAND2XLTS \add_x_22_3/U112  ( .A(\add_x_22_3/n93 ), .B(n1996), .Y(
        \add_x_22_3/n90 ) );
  OR3XLTS U360 ( .A(n2074), .B(\data_cntl/N263 ), .C(n930), .Y(
        \data_cntl/N258 ) );
  NAND2XLTS \add_x_22_5/U112  ( .A(\add_x_22_5/n93 ), .B(n2041), .Y(
        \add_x_22_5/n90 ) );
  NOR2X1TS U392 ( .A(n2585), .B(\data_cntl/N63 ), .Y(\data_cntl/N259 ) );
  NOR3X1TS U393 ( .A(data_to_fft), .B(\data_cntl/N9 ), .C(n2585), .Y(
        \data_cntl/N261 ) );
  NAND3XLTS U395 ( .A(n2071), .B(data_from_fft), .C(data_to_fft), .Y(
        \addr_calc/N216 ) );
  AOI211XLTS U369 ( .A0(n2332), .A1(n935), .B0(n2329), .C0(n1830), .Y(
        \data_cntl/N254 ) );
  CLKINVX1TS U305 ( .A(n899), .Y(n888) );
  CLKINVX2TS U304 ( .A(n870), .Y(n887) );
  NOR3X1TS U378 ( .A(data_to_iir), .B(\data_cntl/N159 ), .C(n932), .Y(
        \data_cntl/N267 ) );
  NOR2X1TS U380 ( .A(\data_cntl/N191 ), .B(n932), .Y(\data_cntl/N265 ) );
  NAND4XLTS U382 ( .A(data_to_iir), .B(data_from_iir), .C(n940), .D(n1830), 
        .Y(\addr_calc/N224 ) );
  CLKAND2X2TS U355 ( .A(n797), .B(fft_put_req_reg), .Y(fft_put_req) );
  OAI211XLTS U302 ( .A0(n888), .A1(n901), .B0(n873), .C0(acc_done), .Y(n890)
         );
  NAND4BXLTS U278 ( .AN(n872), .B(n2055), .C(n2074), .D(n873), .Y(n871) );
  NOR2X1TS U388 ( .A(\data_cntl/N99 ), .B(n1830), .Y(\data_cntl/N262 ) );
  NAND4XLTS U390 ( .A(n2067), .B(data_to_fir), .C(data_from_fir), .D(n2588), 
        .Y(\addr_calc/N220 ) );
  NAND2BXLTS U364 ( .AN(n2323), .B(n2327), .Y(n931) );
  NOR2XLTS U366 ( .A(n2340), .B(n2338), .Y(n933) );
  NAND2BX1TS U370 ( .AN(n2313), .B(n2315), .Y(n935) );
  NOR2XLTS U372 ( .A(n2332), .B(n2329), .Y(n937) );
  AO22X1TS U368 ( .A0(n2332), .A1(n2313), .B0(n2329), .B1(n2315), .Y(n934) );
  NOR2X1TS \add_x_19_4/U38  ( .A(n1929), .B(n2498), .Y(\add_x_19_4/n55 ) );
  NOR3XLTS U375 ( .A(n2334), .B(n2319), .C(n939), .Y(\data_cntl/N251 ) );
  NOR2X1TS \add_x_19_2/U69  ( .A(\add_x_19_2/n81 ), .B(\add_x_19_2/n78 ), .Y(
        \add_x_19_2/n76 ) );
  NAND2XLTS \add_x_22_5/U143  ( .A(\add_x_22_5/n118 ), .B(n2036), .Y(
        \add_x_22_5/n115 ) );
  NAND2X1TS \add_x_19_5/U67  ( .A(\add_x_19_5/n84 ), .B(\add_x_19_5/n76 ), .Y(
        \add_x_19_5/n74 ) );
  NAND2X1TS \add_x_22_1/U7  ( .A(\add_x_22_1/n9 ), .B(n2557), .Y(
        \add_x_22_1/n5 ) );
  NOR2X1TS \add_x_19_3/U34  ( .A(\add_x_19_3/n58 ), .B(\add_x_19_3/n55 ), .Y(
        \add_x_19_3/n53 ) );
  NOR2X1TS \add_x_19_5/U24  ( .A(\add_x_19_5/n51 ), .B(\add_x_19_5/n48 ), .Y(
        \add_x_19_5/n46 ) );
  NAND3XLTS U345 ( .A(n2063), .B(iir_read_done), .C(n924), .Y(n792) );
  NAND2X1TS \add_x_22_2/U123  ( .A(\add_x_22_2/n102 ), .B(n2001), .Y(
        \add_x_22_2/n99 ) );
  NOR2X1TS \add_x_19_1/U24  ( .A(\add_x_19_1/n51 ), .B(\add_x_19_1/n48 ), .Y(
        \add_x_19_1/n46 ) );
  NAND2X1TS \add_x_22_0/U112  ( .A(\add_x_22_0/n93 ), .B(n2049), .Y(
        \add_x_22_0/n90 ) );
  NAND2XLTS U308 ( .A(n870), .B(n884), .Y(n901) );
  NAND2X1TS \add_x_22_1/U81  ( .A(\add_x_22_1/n68 ), .B(n2022), .Y(
        \add_x_22_1/n65 ) );
  NAND2X1TS \add_x_22_1/U59  ( .A(\add_x_22_1/n50 ), .B(
        \addr_calc/fft_write_calc/count[18] ), .Y(\add_x_22_1/n47 ) );
  NAND2X1TS \add_x_22_1/U39  ( .A(\add_x_22_1/n34 ), .B(
        \addr_calc/fft_write_calc/count[22] ), .Y(\add_x_22_1/n31 ) );
  NAND2X1TS \add_x_22_0/U81  ( .A(\add_x_22_0/n68 ), .B(
        \addr_calc/fft_read_calc/count[14] ), .Y(\add_x_22_0/n65 ) );
  CLKAND2X2TS U349 ( .A(n798), .B(fir_put_req_reg), .Y(fir_put_req) );
  NOR2X1TS \add_x_19_1/U178  ( .A(\addr_calc/fft_write_calc/count[10] ), .B(
        n2412), .Y(\add_x_19_1/n144 ) );
  NAND2X1TS \add_x_22_3/U35  ( .A(n1668), .B(n2563), .Y(\add_x_22_3/n28 ) );
  NOR2X1TS \add_x_19_5/U69  ( .A(\add_x_19_5/n81 ), .B(\add_x_19_5/n78 ), .Y(
        \add_x_19_5/n76 ) );
  NAND2X1TS \add_x_19_4/U67  ( .A(\add_x_19_4/n84 ), .B(\add_x_19_4/n76 ), .Y(
        \add_x_19_4/n74 ) );
  NOR2XLTS \add_x_22_2/U132  ( .A(\add_x_22_2/n110 ), .B(\add_x_22_2/n109 ), 
        .Y(\add_x_22_2/n106 ) );
  NAND2XLTS \add_x_22_4/U112  ( .A(\add_x_22_4/n93 ), .B(n2583), .Y(
        \add_x_22_4/n90 ) );
  NAND2XLTS \add_x_22_1/U112  ( .A(\add_x_22_1/n93 ), .B(n2026), .Y(
        \add_x_22_1/n90 ) );
  NAND2XLTS \add_x_22_2/U112  ( .A(\add_x_22_2/n93 ), .B(n1997), .Y(
        \add_x_22_2/n90 ) );
  NAND2XLTS \add_x_22_0/U123  ( .A(\add_x_22_0/n102 ), .B(n2052), .Y(
        \add_x_22_0/n99 ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[6]  ( .D(n996), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[6] ) );
  DFFHQX1TS \addr_calc/iir_write_calc/counter/count_reg[20]  ( .D(n982), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[20] ) );
  DFFHQX1TS \addr_calc/iir_write_calc/counter/count_reg[15]  ( .D(n987), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[15] ) );
  DFFHQX1TS \addr_calc/iir_write_calc/counter/count_reg[16]  ( .D(n986), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[16] ) );
  DFFQX2TS \addr_calc/iir_write_calc/counter/count_reg[29]  ( .D(n973), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[29] ) );
  TBUFX12TS \addr_calc/addr_tri5[21]  ( .A(\addr_calc/iir_read_addr[21] ), 
        .OE(n2769), .Y(addr[21]) );
  TBUFX6TS \addr_calc/addr_tri6[21]  ( .A(\addr_calc/iir_write_addr[21] ), 
        .OE(n2777), .Y(addr[21]) );
  TBUFX6TS \addr_calc/addr_tri4[21]  ( .A(\addr_calc/fir_write_addr[21] ), 
        .OE(n2761), .Y(addr[21]) );
  TBUFX4TS \addr_calc/addr_tri5[24]  ( .A(\addr_calc/iir_read_addr[24] ), .OE(
        n2768), .Y(addr[24]) );
  NAND2X1TS \DP_OP_158_296_6262/U1847  ( .A(\DP_OP_158_296_6262/n1791 ), .B(
        \DP_OP_158_296_6262/n1862 ), .Y(\DP_OP_158_296_6262/n1861 ) );
  NAND2X1TS \add_x_19_4/U26  ( .A(\add_x_19_4/n195 ), .B(\add_x_19_4/n49 ), 
        .Y(\add_x_19_4/n4 ) );
  NAND2X1TS \add_x_19_4/U50  ( .A(\add_x_19_4/n198 ), .B(\add_x_19_4/n64 ), 
        .Y(\add_x_19_4/n7 ) );
  OAI21X1TS \add_x_19_4/U136  ( .A0(\add_x_19_4/n120 ), .A1(\add_x_19_4/n124 ), 
        .B0(\add_x_19_4/n121 ), .Y(\add_x_19_4/n119 ) );
  NAND2X1TS \add_x_19_4/U22  ( .A(\add_x_19_4/n72 ), .B(\add_x_19_4/n46 ), .Y(
        \add_x_19_4/n44 ) );
  OAI21X1TS \add_x_19_4/U25  ( .A0(\add_x_19_4/n52 ), .A1(\add_x_19_4/n48 ), 
        .B0(\add_x_19_4/n49 ), .Y(\add_x_19_4/n47 ) );
  XNOR2X1TS \add_x_19_4/U128  ( .A(\add_x_19_4/n122 ), .B(\add_x_19_4/n17 ), 
        .Y(\addr_calc/iir_read_addr[15] ) );
  OAI21X1TS \add_x_19_4/U142  ( .A0(\add_x_19_4/n125 ), .A1(\add_x_19_4/n123 ), 
        .B0(\add_x_19_4/n124 ), .Y(\add_x_19_4/n122 ) );
  NAND2X1TS \add_x_19_4/U137  ( .A(\add_x_19_4/n208 ), .B(\add_x_19_4/n121 ), 
        .Y(\add_x_19_4/n17 ) );
  NOR2X1TS \add_x_22_1/U132  ( .A(\add_x_22_1/n110 ), .B(\add_x_22_1/n109 ), 
        .Y(\add_x_22_1/n106 ) );
  NOR2X1TS \DP_OP_159_297_3515/U941  ( .A(\DP_OP_159_297_3515/n957 ), .B(
        \DP_OP_159_297_3515/n943 ), .Y(\DP_OP_159_297_3515/n942 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1874  ( .A(\DP_OP_158_296_6262/n1883 ), .B(
        \DP_OP_158_296_6262/n1904 ), .Y(\DP_OP_158_296_6262/n1882 ) );
  AOI21X1TS \add_x_19_0/U134  ( .A0(\add_x_19_0/n118 ), .A1(\add_x_19_0/n127 ), 
        .B0(\add_x_19_0/n119 ), .Y(\add_x_19_0/n117 ) );
  OAI21X1TS \add_x_19_0/U136  ( .A0(\add_x_19_0/n120 ), .A1(\add_x_19_0/n124 ), 
        .B0(\add_x_19_0/n121 ), .Y(\add_x_19_0/n119 ) );
  OAI21X1TS \add_x_19_0/U202  ( .A0(\add_x_19_0/n162 ), .A1(\add_x_19_0/n166 ), 
        .B0(\add_x_19_0/n163 ), .Y(\add_x_19_0/n161 ) );
  NAND2X2TS \DP_OP_158_296_6262/U1090  ( .A(\DP_OP_158_296_6262/n1073 ), .B(
        \DP_OP_158_296_6262/n1174 ), .Y(\DP_OP_158_296_6262/n1071 ) );
  NOR2X2TS \DP_OP_158_296_6262/U1092  ( .A(\DP_OP_158_296_6262/n1075 ), .B(
        \DP_OP_158_296_6262/n1132 ), .Y(\DP_OP_158_296_6262/n1073 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U906  ( .A(n1778), .B(
        \addr_calc/fft_read_calc/count[31] ), .Y(\DP_OP_158_296_6262/n899 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1185  ( .A(n1659), .B(
        \addr_calc/fft_read_calc/count[13] ), .Y(\DP_OP_158_296_6262/n1160 )
         );
  XNOR2X1TS \DP_OP_158_296_6262/U1219  ( .A(n1656), .B(n1972), .Y(
        \DP_OP_158_296_6262/n1191 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1229  ( .A(n1469), .B(n2560), .Y(
        \DP_OP_158_296_6262/n1200 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1239  ( .A(n2598), .B(n2049), .Y(
        \DP_OP_158_296_6262/n1209 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1255  ( .A(n1602), .B(n1599), .Y(
        \DP_OP_158_296_6262/n1223 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1277  ( .A(n1600), .B(n1601), .Y(
        \DP_OP_158_296_6262/n1243 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1295  ( .A(\DP_OP_158_296_6262/n1265 ), .B(
        n1598), .Y(\DP_OP_158_296_6262/n1259 ) );
  NOR2X1TS \DP_OP_158_296_6262/U1302  ( .A(\DP_OP_158_296_6262/n1267 ), .B(
        \DP_OP_158_296_6262/n1269 ), .Y(\DP_OP_158_296_6262/n1265 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1304  ( .A(\addr_calc/fft_read_calc/count[1] ), .B(n2597), .Y(\DP_OP_158_296_6262/n1267 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1311  ( .A(n2372), .B(n2058), .Y(
        \DP_OP_158_296_6262/n1269 ) );
  NOR2X1TS \DP_OP_158_296_6262/U1821  ( .A(\DP_OP_158_296_6262/n1792 ), .B(
        n1807), .Y(\DP_OP_158_296_6262/n1842 ) );
  NAND2X1TS \add_x_19_3/U71  ( .A(\add_x_19_3/n200 ), .B(\add_x_19_3/n79 ), 
        .Y(\add_x_19_3/n9 ) );
  AOI21X1TS \add_x_19_3/U82  ( .A0(\add_x_19_3/n92 ), .A1(\add_x_19_3/n84 ), 
        .B0(\add_x_19_3/n85 ), .Y(\add_x_19_3/n83 ) );
  OAI21X1TS \add_x_19_3/U97  ( .A0(\add_x_19_3/n113 ), .A1(\add_x_19_3/n93 ), 
        .B0(\add_x_19_3/n94 ), .Y(\add_x_19_3/n92 ) );
  NAND2X1TS \add_x_19_5/U2  ( .A(n1590), .B(\add_x_19_5/n34 ), .Y(
        \add_x_19_5/n1 ) );
  NAND2XLTS \add_x_19_5/U5  ( .A(n1857), .B(n2382), .Y(\add_x_19_5/n34 ) );
  OAI21X2TS \add_x_19_4/U198  ( .A0(\add_x_19_4/n178 ), .A1(\add_x_19_4/n158 ), 
        .B0(\add_x_19_4/n159 ), .Y(\add_x_19_4/n157 ) );
  NAND2X1TS \add_x_19_4/U199  ( .A(\add_x_19_4/n168 ), .B(\add_x_19_4/n160 ), 
        .Y(\add_x_19_4/n158 ) );
  AOI21X1TS \add_x_19_4/U200  ( .A0(\add_x_19_4/n160 ), .A1(\add_x_19_4/n169 ), 
        .B0(\add_x_19_4/n161 ), .Y(\add_x_19_4/n159 ) );
  OAI21X1TS \add_x_19_4/U202  ( .A0(\add_x_19_4/n162 ), .A1(\add_x_19_4/n166 ), 
        .B0(\add_x_19_4/n163 ), .Y(\add_x_19_4/n161 ) );
  OAI21X1TS \add_x_19_4/U216  ( .A0(\add_x_19_4/n170 ), .A1(\add_x_19_4/n176 ), 
        .B0(\add_x_19_4/n171 ), .Y(\add_x_19_4/n169 ) );
  OAI21X1TS \add_x_19_5/U76  ( .A0(\add_x_19_5/n83 ), .A1(\add_x_19_5/n81 ), 
        .B0(\add_x_19_5/n82 ), .Y(\add_x_19_5/n80 ) );
  NAND2X1TS \add_x_19_5/U71  ( .A(\add_x_19_5/n200 ), .B(\add_x_19_5/n79 ), 
        .Y(\add_x_19_5/n9 ) );
  AOI21X1TS \add_x_19_3/U165  ( .A0(\add_x_19_3/n137 ), .A1(\add_x_19_3/n150 ), 
        .B0(\add_x_19_3/n138 ), .Y(\add_x_19_3/n136 ) );
  OAI21X1TS \add_x_19_3/U167  ( .A0(\add_x_19_3/n139 ), .A1(\add_x_19_3/n145 ), 
        .B0(\add_x_19_3/n140 ), .Y(\add_x_19_3/n138 ) );
  XOR2X1TS \add_x_22_5/U42  ( .A(\add_x_22_5/n38 ), .B(n1961), .Y(
        \addr_calc/iir_write_calc/counter/N64 ) );
  NAND2X1TS \add_x_22_5/U48  ( .A(\add_x_22_5/n41 ), .B(
        \addr_calc/iir_write_calc/count[20] ), .Y(\add_x_22_5/n38 ) );
  NOR2X1TS \DP_OP_159_297_3515/U881  ( .A(n2551), .B(\DP_OP_159_297_3515/n901 ), .Y(\DP_OP_159_297_3515/n900 ) );
  NOR2X1TS \DP_OP_159_297_3515/U883  ( .A(\DP_OP_159_297_3515/n915 ), .B(
        \DP_OP_159_297_3515/n903 ), .Y(\DP_OP_159_297_3515/n902 ) );
  NAND2X1TS \DP_OP_159_297_3515/U884  ( .A(n1562), .B(n1807), .Y(
        \DP_OP_159_297_3515/n903 ) );
  NAND2X1TS \DP_OP_159_297_3515/U904  ( .A(n1485), .B(n1664), .Y(
        \DP_OP_159_297_3515/n915 ) );
  OAI21X2TS \add_x_19_3/U198  ( .A0(\add_x_19_3/n178 ), .A1(\add_x_19_3/n158 ), 
        .B0(\add_x_19_3/n159 ), .Y(\add_x_19_3/n157 ) );
  NAND2X1TS \add_x_19_3/U199  ( .A(\add_x_19_3/n168 ), .B(\add_x_19_3/n160 ), 
        .Y(\add_x_19_3/n158 ) );
  AOI21X1TS \add_x_19_3/U200  ( .A0(\add_x_19_3/n160 ), .A1(\add_x_19_3/n169 ), 
        .B0(\add_x_19_3/n161 ), .Y(\add_x_19_3/n159 ) );
  OAI21X1TS \add_x_19_3/U202  ( .A0(\add_x_19_3/n162 ), .A1(\add_x_19_3/n166 ), 
        .B0(\add_x_19_3/n163 ), .Y(\add_x_19_3/n161 ) );
  NOR2X1TS \add_x_19_3/U201  ( .A(\add_x_19_3/n165 ), .B(\add_x_19_3/n162 ), 
        .Y(\add_x_19_3/n160 ) );
  NAND2X1TS \add_x_19_2/U2  ( .A(n1560), .B(\add_x_19_2/n34 ), .Y(
        \add_x_19_2/n1 ) );
  NAND2XLTS \add_x_19_2/U5  ( .A(n2549), .B(n2380), .Y(\add_x_19_2/n34 ) );
  AOI21X1TS \add_x_19_0/U82  ( .A0(\add_x_19_0/n92 ), .A1(\add_x_19_0/n84 ), 
        .B0(\add_x_19_0/n85 ), .Y(\add_x_19_0/n83 ) );
  OAI21X1TS \add_x_19_0/U97  ( .A0(\add_x_19_0/n113 ), .A1(\add_x_19_0/n93 ), 
        .B0(\add_x_19_0/n94 ), .Y(\add_x_19_0/n92 ) );
  OAI21X2TS \add_x_19_0/U198  ( .A0(\add_x_19_0/n178 ), .A1(\add_x_19_0/n158 ), 
        .B0(\add_x_19_0/n159 ), .Y(\add_x_19_0/n157 ) );
  XNOR2X1TS \add_x_19_5/U95  ( .A(\add_x_19_5/n99 ), .B(\add_x_19_5/n13 ), .Y(
        \addr_calc/iir_write_addr[19] ) );
  OAI21X1TS \add_x_19_5/U107  ( .A0(\add_x_19_5/n102 ), .A1(\add_x_19_5/n100 ), 
        .B0(\add_x_19_5/n101 ), .Y(\add_x_19_5/n99 ) );
  NAND2X1TS \add_x_19_5/U102  ( .A(\add_x_19_5/n204 ), .B(\add_x_19_5/n98 ), 
        .Y(\add_x_19_5/n13 ) );
  NAND2X1TS \add_x_19_1/U36  ( .A(\add_x_19_1/n196 ), .B(\add_x_19_1/n56 ), 
        .Y(\add_x_19_1/n5 ) );
  NOR2X1TS \add_x_19_1/U232  ( .A(\add_x_19_1/n184 ), .B(\add_x_19_1/n181 ), 
        .Y(\add_x_19_1/n179 ) );
  OAI21X1TS \add_x_19_1/U233  ( .A0(\add_x_19_1/n181 ), .A1(\add_x_19_1/n185 ), 
        .B0(\add_x_19_1/n182 ), .Y(\add_x_19_1/n180 ) );
  OAI21X1TS \add_x_19_0/U150  ( .A0(\add_x_19_0/n128 ), .A1(\add_x_19_0/n132 ), 
        .B0(\add_x_19_0/n129 ), .Y(\add_x_19_0/n127 ) );
  NOR2X1TS \add_x_19_3/U232  ( .A(\add_x_19_3/n184 ), .B(\add_x_19_3/n181 ), 
        .Y(\add_x_19_3/n179 ) );
  OAI21X1TS \add_x_19_3/U233  ( .A0(\add_x_19_3/n181 ), .A1(\add_x_19_3/n185 ), 
        .B0(\add_x_19_3/n182 ), .Y(\add_x_19_3/n180 ) );
  NOR2X1TS \add_x_19_1/U215  ( .A(\add_x_19_1/n175 ), .B(\add_x_19_1/n170 ), 
        .Y(\add_x_19_1/n168 ) );
  AOI21X1TS \add_x_19_0/U47  ( .A0(\add_x_19_0/n69 ), .A1(\add_x_19_0/n61 ), 
        .B0(\add_x_19_0/n62 ), .Y(\add_x_19_0/n60 ) );
  NOR2X1TS \add_x_19_0/U65  ( .A(\add_x_19_0/n93 ), .B(\add_x_19_0/n74 ), .Y(
        \add_x_19_0/n72 ) );
  NAND2X1TS \add_x_19_0/U67  ( .A(\add_x_19_0/n84 ), .B(\add_x_19_0/n76 ), .Y(
        \add_x_19_0/n74 ) );
  OAI21X1TS \add_x_19_0/U66  ( .A0(\add_x_19_0/n94 ), .A1(\add_x_19_0/n74 ), 
        .B0(\add_x_19_0/n75 ), .Y(\add_x_19_0/n73 ) );
  AOI21X1TS \add_x_19_0/U68  ( .A0(\add_x_19_0/n85 ), .A1(\add_x_19_0/n76 ), 
        .B0(\add_x_19_0/n77 ), .Y(\add_x_19_0/n75 ) );
  OAI21X1TS \add_x_19_0/U70  ( .A0(\add_x_19_0/n78 ), .A1(\add_x_19_0/n82 ), 
        .B0(\add_x_19_0/n79 ), .Y(\add_x_19_0/n77 ) );
  NAND2X1TS \add_x_19_2/U22  ( .A(\add_x_19_2/n72 ), .B(\add_x_19_2/n46 ), .Y(
        \add_x_19_2/n44 ) );
  OAI21X1TS \add_x_19_2/U25  ( .A0(\add_x_19_2/n52 ), .A1(\add_x_19_2/n48 ), 
        .B0(\add_x_19_2/n49 ), .Y(\add_x_19_2/n47 ) );
  NOR2X1TS \add_x_19_4/U232  ( .A(\add_x_19_4/n184 ), .B(\add_x_19_4/n181 ), 
        .Y(\add_x_19_4/n179 ) );
  OAI21X1TS \add_x_19_4/U233  ( .A0(\add_x_19_4/n181 ), .A1(\add_x_19_4/n185 ), 
        .B0(\add_x_19_4/n182 ), .Y(\add_x_19_4/n180 ) );
  NOR2X1TS \add_x_19_0/U135  ( .A(\add_x_19_0/n123 ), .B(\add_x_19_0/n120 ), 
        .Y(\add_x_19_0/n118 ) );
  NOR2X1TS \add_x_19_1/U166  ( .A(\add_x_19_1/n144 ), .B(\add_x_19_1/n139 ), 
        .Y(\add_x_19_1/n137 ) );
  AOI21X1TS \add_x_19_2/U165  ( .A0(\add_x_19_2/n137 ), .A1(\add_x_19_2/n150 ), 
        .B0(\add_x_19_2/n138 ), .Y(\add_x_19_2/n136 ) );
  OAI21X1TS \add_x_19_2/U167  ( .A0(\add_x_19_2/n139 ), .A1(\add_x_19_2/n145 ), 
        .B0(\add_x_19_2/n140 ), .Y(\add_x_19_2/n138 ) );
  NOR2X1TS \add_x_19_1/U135  ( .A(\add_x_19_1/n123 ), .B(\add_x_19_1/n120 ), 
        .Y(\add_x_19_1/n118 ) );
  NOR2X1TS \add_x_19_2/U24  ( .A(\add_x_19_2/n51 ), .B(\add_x_19_2/n48 ), .Y(
        \add_x_19_2/n46 ) );
  NOR2X1TS \add_x_19_1/U201  ( .A(\add_x_19_1/n165 ), .B(\add_x_19_1/n162 ), 
        .Y(\add_x_19_1/n160 ) );
  OAI21X1TS \add_x_19_2/U216  ( .A0(\add_x_19_2/n170 ), .A1(\add_x_19_2/n176 ), 
        .B0(\add_x_19_2/n171 ), .Y(\add_x_19_2/n169 ) );
  NOR2X1TS \add_x_19_2/U219  ( .A(n1904), .B(n2484), .Y(\add_x_19_2/n170 ) );
  OAI21X1TS \add_x_19_2/U66  ( .A0(\add_x_19_2/n94 ), .A1(\add_x_19_2/n74 ), 
        .B0(\add_x_19_2/n75 ), .Y(\add_x_19_2/n73 ) );
  AOI21X1TS \add_x_19_2/U68  ( .A0(\add_x_19_2/n76 ), .A1(\add_x_19_2/n85 ), 
        .B0(\add_x_19_2/n77 ), .Y(\add_x_19_2/n75 ) );
  OAI21X1TS \add_x_19_2/U70  ( .A0(\add_x_19_2/n78 ), .A1(\add_x_19_2/n82 ), 
        .B0(\add_x_19_2/n79 ), .Y(\add_x_19_2/n77 ) );
  OAI21X1TS \add_x_19_2/U84  ( .A0(\add_x_19_2/n86 ), .A1(\add_x_19_2/n90 ), 
        .B0(\add_x_19_2/n87 ), .Y(\add_x_19_2/n85 ) );
  AOI21X1TS \add_x_19_5/U148  ( .A0(\add_x_19_5/n134 ), .A1(\add_x_19_5/n126 ), 
        .B0(\add_x_19_5/n127 ), .Y(\add_x_19_5/n125 ) );
  OAI21X1TS \add_x_19_5/U25  ( .A0(\add_x_19_5/n52 ), .A1(\add_x_19_5/n48 ), 
        .B0(\add_x_19_5/n49 ), .Y(\add_x_19_5/n47 ) );
  AOI21X1TS \add_x_19_5/U68  ( .A0(\add_x_19_5/n76 ), .A1(\add_x_19_5/n85 ), 
        .B0(\add_x_19_5/n77 ), .Y(\add_x_19_5/n75 ) );
  OAI21X1TS \add_x_19_5/U70  ( .A0(\add_x_19_5/n78 ), .A1(\add_x_19_5/n82 ), 
        .B0(\add_x_19_5/n79 ), .Y(\add_x_19_5/n77 ) );
  OAI21X1TS \add_x_19_5/U84  ( .A0(\add_x_19_5/n86 ), .A1(\add_x_19_5/n90 ), 
        .B0(\add_x_19_5/n87 ), .Y(\add_x_19_5/n85 ) );
  NAND2X1TS \add_x_19_1/U71  ( .A(\add_x_19_1/n200 ), .B(\add_x_19_1/n79 ), 
        .Y(\add_x_19_1/n9 ) );
  DFFTRX2TS \addr_calc/fft_write_calc/counter/done_reg  ( .D(n1675), .RN(n2072), .CK(clk), .Q(n1478), .QN(n1828) );
  DFFTRX2TS \addr_calc/iir_read_calc/counter/done_reg  ( .D(n1781), .RN(n2063), 
        .CK(clk), .Q(iir_read_done), .QN(n898) );
  DFFXLTS \pla_top/fft_enable_reg  ( .D(n1131), .CK(clk), .Q(fft_enable), .QN(
        n2070) );
  DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[14]  ( .D(n957), .CK(clk), .Q(\addr_calc/iir_read_calc/count[14] ) );
  TBUFX4TS \addr_calc/addr_tri[22]  ( .A(\addr_calc/fft_read_addr[22] ), .OE(
        n2737), .Y(addr[22]) );
  TBUFX4TS \addr_calc/addr_tri6[22]  ( .A(\addr_calc/iir_write_addr[22] ), 
        .OE(n2777), .Y(addr[22]) );
  DFFQX4TS \addr_calc/fir_read_calc/counter/count_reg[7]  ( .D(n1091), .CK(clk), .Q(\addr_calc/fir_read_calc/count[7] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[31]  ( .D(n1035), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[31] ) );
  DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[23]  ( .D(n1011), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[23] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[23]  ( .D(n979), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[23] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[24]  ( .D(n978), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[24] ) );
  TBUFX12TS \addr_calc/addr_tri5[19]  ( .A(\addr_calc/iir_read_addr[19] ), 
        .OE(n2770), .Y(addr[19]) );
  TBUFX6TS \addr_calc/addr_tri6[19]  ( .A(\addr_calc/iir_write_addr[19] ), 
        .OE(n2778), .Y(addr[19]) );
  TBUFX6TS \addr_calc/addr_tri4[19]  ( .A(\addr_calc/fir_write_addr[19] ), 
        .OE(n2762), .Y(addr[19]) );
  TBUFX4TS \addr_calc/addr_tri3[18]  ( .A(\addr_calc/fir_read_addr[18] ), .OE(
        n2754), .Y(addr[18]) );
  DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[17]  ( .D(n954), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[17] ) );
  TBUFX4TS \addr_calc/addr_tri6[18]  ( .A(\addr_calc/iir_write_addr[18] ), 
        .OE(n2778), .Y(addr[18]) );
  TBUFX4TS \addr_calc/addr_tri2[18]  ( .A(\addr_calc/fft_write_addr[18] ), 
        .OE(n2746), .Y(addr[18]) );
  TBUFX4TS \addr_calc/addr_tri4[13]  ( .A(\addr_calc/fir_write_addr[13] ), 
        .OE(n2763), .Y(addr[13]) );
  TBUFX4TS \addr_calc/addr_tri2[13]  ( .A(\addr_calc/fft_write_addr[13] ), 
        .OE(n2747), .Y(addr[13]) );
  TBUFX6TS \addr_calc/addr_tri2[30]  ( .A(\addr_calc/fft_write_addr[30] ), 
        .OE(n2743), .Y(addr[30]) );
  DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[23]  ( .D(n948), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[23] ) );
  DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[15]  ( .D(n956), .CK(clk), .Q(\addr_calc/iir_read_calc/count[15] ) );
  TBUFX12TS \addr_calc/addr_tri5[25]  ( .A(\addr_calc/iir_read_addr[25] ), 
        .OE(n2768), .Y(addr[25]) );
  TBUFX6TS \addr_calc/addr_tri[25]  ( .A(\addr_calc/fft_read_addr[25] ), .OE(
        n2736), .Y(addr[25]) );
  TBUFX6TS \addr_calc/addr_tri[28]  ( .A(\addr_calc/fft_read_addr[28] ), .OE(
        n2735), .Y(addr[28]) );
  TBUFX12TS \addr_calc/addr_tri5[28]  ( .A(\addr_calc/iir_read_addr[28] ), 
        .OE(n2767), .Y(addr[28]) );
  TBUFX12TS \addr_calc/addr_tri2[28]  ( .A(\addr_calc/fft_write_addr[28] ), 
        .OE(n2743), .Y(addr[28]) );
  TBUFX4TS \addr_calc/addr_tri2[14]  ( .A(\addr_calc/fft_write_addr[14] ), 
        .OE(n2747), .Y(addr[14]) );
  TBUFX4TS \addr_calc/addr_tri2[17]  ( .A(\addr_calc/fft_write_addr[17] ), 
        .OE(n2746), .Y(addr[17]) );
  TBUFX6TS \addr_calc/addr_tri2[26]  ( .A(\addr_calc/fft_write_addr[26] ), 
        .OE(n2744), .Y(addr[26]) );
  TBUFX12TS \addr_calc/addr_tri2[15]  ( .A(\addr_calc/fft_write_addr[15] ), 
        .OE(n2747), .Y(addr[15]) );
  DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[22]  ( .D(n949), .CK(
        clk), .Q(\addr_calc/iir_read_calc/count[22] ) );
  TBUFX12TS \addr_calc/addr_tri3[21]  ( .A(\addr_calc/fir_read_addr[21] ), 
        .OE(n2753), .Y(addr[21]) );
  TBUFX2TS \addr_calc/addr_tri[14]  ( .A(\addr_calc/fft_read_addr[14] ), .OE(
        n2739), .Y(addr[14]) );
  TBUFX4TS \addr_calc/addr_tri6[30]  ( .A(\addr_calc/iir_write_addr[30] ), 
        .OE(n2775), .Y(addr[30]) );
  TBUFX8TS \addr_calc/addr_tri4[27]  ( .A(\addr_calc/fir_write_addr[27] ), 
        .OE(n2760), .Y(addr[27]) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[2]  ( .D(n1000), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[2] ) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[13]  ( .D(n989), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[13] ) );
  TBUFX4TS \addr_calc/addr_tri5[17]  ( .A(\addr_calc/iir_read_addr[17] ), .OE(
        n2770), .Y(addr[17]) );
  TBUFX6TS \addr_calc/addr_tri5[22]  ( .A(\addr_calc/iir_read_addr[22] ), .OE(
        n2769), .Y(addr[22]) );
  TBUFX4TS \addr_calc/addr_tri3[22]  ( .A(\addr_calc/fir_read_addr[22] ), .OE(
        n2753), .Y(addr[22]) );
  TBUFX12TS \addr_calc/addr_tri2[21]  ( .A(\addr_calc/fft_write_addr[21] ), 
        .OE(n2745), .Y(addr[21]) );
  TBUFX2TS \addr_calc/addr_tri[18]  ( .A(\addr_calc/fft_read_addr[18] ), .OE(
        n2738), .Y(addr[18]) );
  TBUFX2TS \addr_calc/addr_tri4[18]  ( .A(\addr_calc/fir_write_addr[18] ), 
        .OE(n2762), .Y(addr[18]) );
  TBUFX12TS \addr_calc/addr_tri[23]  ( .A(\addr_calc/fft_read_addr[23] ), .OE(
        n2737), .Y(addr[23]) );
  TBUFX12TS \addr_calc/addr_tri3[23]  ( .A(\addr_calc/fir_read_addr[23] ), 
        .OE(n2753), .Y(addr[23]) );
  TBUFX12TS \addr_calc/addr_tri6[23]  ( .A(\addr_calc/iir_write_addr[23] ), 
        .OE(n2777), .Y(addr[23]) );
  XOR2X1TS \add_x_22_4/U42  ( .A(\add_x_22_4/n38 ), .B(n1923), .Y(
        \addr_calc/iir_read_calc/counter/N64 ) );
  NAND2X1TS \add_x_22_4/U48  ( .A(\add_x_22_4/n41 ), .B(
        \addr_calc/iir_read_calc/count[20] ), .Y(\add_x_22_4/n38 ) );
  XNOR2X1TS \DP_OP_159_297_3515/U341  ( .A(n2609), .B(
        \addr_calc/iir_read_calc/count[7] ), .Y(\DP_OP_159_297_3515/n312 ) );
  NAND2X1TS \DP_OP_159_297_3515/U347  ( .A(n1247), .B(n1249), .Y(
        \DP_OP_159_297_3515/n317 ) );
  NAND2X1TS \DP_OP_159_297_3515/U377  ( .A(\DP_OP_159_297_3515/n349 ), .B(
        n1246), .Y(\DP_OP_159_297_3515/n343 ) );
  XNOR2X1TS \DP_OP_159_297_3515/U374  ( .A(n2611), .B(n1902), .Y(
        \DP_OP_159_297_3515/n341 ) );
  NOR2X1TS \DP_OP_159_297_3515/U384  ( .A(\DP_OP_159_297_3515/n351 ), .B(
        \DP_OP_159_297_3515/n353 ), .Y(\DP_OP_159_297_3515/n349 ) );
  XNOR2X1TS \DP_OP_159_297_3515/U386  ( .A(n2374), .B(
        \addr_calc/iir_read_calc/count[1] ), .Y(\DP_OP_159_297_3515/n351 ) );
  NAND2X1TS \DP_OP_159_297_3515/U1003  ( .A(n1520), .B(n1529), .Y(
        \DP_OP_159_297_3515/n986 ) );
  XOR2X1TS \add_x_22_3/U115  ( .A(\add_x_22_3/n99 ), .B(\add_x_22_3/n98 ), .Y(
        \addr_calc/fir_write_calc/counter/N50 ) );
  NAND2XLTS \add_x_22_3/U123  ( .A(\add_x_22_3/n102 ), .B(n1993), .Y(
        \add_x_22_3/n99 ) );
  XOR2X1TS \add_x_22_3/U100  ( .A(\add_x_22_3/n85 ), .B(\add_x_22_3/n84 ), .Y(
        \addr_calc/fir_write_calc/counter/N53 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1354  ( .A(n1778), .B(
        \addr_calc/fir_write_calc/count[31] ), .Y(\DP_OP_158_296_6262/n1346 )
         );
  NOR2X1TS \DP_OP_158_296_6262/U1723  ( .A(\DP_OP_158_296_6262/n1690 ), .B(
        \DP_OP_158_296_6262/n1706 ), .Y(\DP_OP_158_296_6262/n1688 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1406  ( .A(n1775), .B(
        \addr_calc/fir_write_calc/count[28] ), .Y(\DP_OP_158_296_6262/n1395 )
         );
  XNOR2X1TS \DP_OP_158_296_6262/U1594  ( .A(n2594), .B(n2564), .Y(
        \DP_OP_158_296_6262/n1571 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1621  ( .A(n1657), .B(n2003), .Y(
        \DP_OP_158_296_6262/n1596 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1607  ( .A(n1658), .B(
        \addr_calc/fir_write_calc/count[15] ), .Y(\DP_OP_158_296_6262/n1583 )
         );
  XNOR2X1TS \DP_OP_158_296_6262/U1655  ( .A(n1660), .B(n1877), .Y(
        \DP_OP_158_296_6262/n1627 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1687  ( .A(n2598), .B(n1996), .Y(
        \DP_OP_158_296_6262/n1656 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1695  ( .A(n1651), .B(n1869), .Y(
        \DP_OP_158_296_6262/n1663 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1703  ( .A(n1239), .B(n1236), .Y(
        \DP_OP_158_296_6262/n1670 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1725  ( .A(n1237), .B(n1238), .Y(
        \DP_OP_158_296_6262/n1690 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1743  ( .A(\DP_OP_158_296_6262/n1712 ), .B(
        n1235), .Y(\DP_OP_158_296_6262/n1706 ) );
  NOR2X1TS \DP_OP_158_296_6262/U1750  ( .A(\DP_OP_158_296_6262/n1714 ), .B(
        \DP_OP_158_296_6262/n1716 ), .Y(\DP_OP_158_296_6262/n1712 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U1752  ( .A(n2597), .B(n1868), .Y(
        \DP_OP_158_296_6262/n1714 ) );
  NOR2X8TS \DP_OP_158_296_6262/U2008  ( .A(\DP_OP_158_296_6262/n2011 ), .B(
        \DP_OP_158_296_6262/n1987 ), .Y(\DP_OP_158_296_6262/n1986 ) );
  XNOR2X1TS \add_x_22_1/U58  ( .A(\add_x_22_1/n50 ), .B(n2019), .Y(
        \addr_calc/fft_write_calc/counter/N61 ) );
  NOR2X2TS \DP_OP_158_296_6262/U644  ( .A(\DP_OP_158_296_6262/n628 ), .B(
        \DP_OP_158_296_6262/n685 ), .Y(\DP_OP_158_296_6262/n626 ) );
  NOR2X2TS \DP_OP_158_296_6262/U753  ( .A(\DP_OP_158_296_6262/n729 ), .B(
        \DP_OP_158_296_6262/n765 ), .Y(\DP_OP_158_296_6262/n727 ) );
  NAND2X1TS \DP_OP_158_296_6262/U795  ( .A(\DP_OP_158_296_6262/n767 ), .B(
        \DP_OP_158_296_6262/n794 ), .Y(\DP_OP_158_296_6262/n765 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U458  ( .A(n1778), .B(
        \addr_calc/fft_write_calc/count[31] ), .Y(\DP_OP_158_296_6262/n452 )
         );
  NOR2X1TS \DP_OP_158_296_6262/U827  ( .A(\DP_OP_158_296_6262/n796 ), .B(
        \DP_OP_158_296_6262/n812 ), .Y(\DP_OP_158_296_6262/n794 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U698  ( .A(n2594), .B(n2567), .Y(
        \DP_OP_158_296_6262/n677 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U737  ( .A(n1927), .B(n1659), .Y(
        \DP_OP_158_296_6262/n713 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U771  ( .A(n1656), .B(n1932), .Y(
        \DP_OP_158_296_6262/n744 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U781  ( .A(n1469), .B(n1934), .Y(
        \DP_OP_158_296_6262/n753 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U791  ( .A(n2598), .B(n2026), .Y(
        \DP_OP_158_296_6262/n762 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U799  ( .A(n1651), .B(n1936), .Y(
        \DP_OP_158_296_6262/n769 ) );
  NAND2X1TS \DP_OP_158_296_6262/U807  ( .A(n1212), .B(n1209), .Y(
        \DP_OP_158_296_6262/n776 ) );
  NAND2X1TS \DP_OP_158_296_6262/U829  ( .A(n1210), .B(n1211), .Y(
        \DP_OP_158_296_6262/n796 ) );
  NAND2X1TS \DP_OP_158_296_6262/U847  ( .A(\DP_OP_158_296_6262/n818 ), .B(
        n1208), .Y(\DP_OP_158_296_6262/n812 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U510  ( .A(n1775), .B(
        \addr_calc/fft_write_calc/count[28] ), .Y(\DP_OP_158_296_6262/n501 )
         );
  NOR2X1TS \DP_OP_158_296_6262/U854  ( .A(\DP_OP_158_296_6262/n820 ), .B(
        \DP_OP_158_296_6262/n822 ), .Y(\DP_OP_158_296_6262/n818 ) );
  XNOR2X1TS \DP_OP_158_296_6262/U856  ( .A(n2597), .B(n1941), .Y(
        \DP_OP_158_296_6262/n820 ) );
  NAND2X1TS \DP_OP_158_296_6262/U1883  ( .A(\DP_OP_158_296_6262/n1904 ), .B(
        \DP_OP_158_296_6262/n1890 ), .Y(\DP_OP_158_296_6262/n1889 ) );
  XOR2X1TS \add_x_22_4/U131  ( .A(\add_x_22_4/n110 ), .B(\add_x_22_4/n109 ), 
        .Y(\addr_calc/iir_read_calc/counter/N47 ) );
  XNOR2X1TS \add_x_22_4/U122  ( .A(\add_x_22_4/n102 ), .B(\add_x_22_4/n101 ), 
        .Y(\addr_calc/iir_read_calc/counter/N49 ) );
  XOR2X1TS \add_x_22_3/U72  ( .A(\add_x_22_3/n65 ), .B(n1882), .Y(
        \addr_calc/fir_write_calc/counter/N58 ) );
  OAI21X1TS \add_x_19_2/U31  ( .A0(\add_x_19_2/n68 ), .A1(\add_x_19_2/n51 ), 
        .B0(\add_x_19_2/n52 ), .Y(\add_x_19_2/n50 ) );
  NAND2X1TS \add_x_19_2/U26  ( .A(\add_x_19_2/n195 ), .B(\add_x_19_2/n49 ), 
        .Y(\add_x_19_2/n4 ) );
  OAI21X1TS \add_x_19_2/U55  ( .A0(\add_x_19_2/n68 ), .A1(\add_x_19_2/n66 ), 
        .B0(\add_x_19_2/n67 ), .Y(\add_x_19_2/n65 ) );
  NAND2X1TS \add_x_19_2/U50  ( .A(\add_x_19_2/n198 ), .B(\add_x_19_2/n64 ), 
        .Y(\add_x_19_2/n7 ) );
  NOR2X1TS \add_x_19_2/U131  ( .A(\add_x_19_2/n135 ), .B(\add_x_19_2/n116 ), 
        .Y(\add_x_19_2/n114 ) );
  AOI21X1TS \add_x_19_2/U134  ( .A0(\add_x_19_2/n118 ), .A1(\add_x_19_2/n127 ), 
        .B0(\add_x_19_2/n119 ), .Y(\add_x_19_2/n117 ) );
  OAI21X1TS \add_x_19_2/U136  ( .A0(\add_x_19_2/n120 ), .A1(\add_x_19_2/n124 ), 
        .B0(\add_x_19_2/n121 ), .Y(\add_x_19_2/n119 ) );
  OAI21X2TS \add_x_19_2/U198  ( .A0(\add_x_19_2/n178 ), .A1(\add_x_19_2/n158 ), 
        .B0(\add_x_19_2/n159 ), .Y(\add_x_19_2/n157 ) );
  AOI21X1TS \add_x_19_2/U200  ( .A0(\add_x_19_2/n160 ), .A1(\add_x_19_2/n169 ), 
        .B0(\add_x_19_2/n161 ), .Y(\add_x_19_2/n159 ) );
  OAI21X1TS \add_x_19_2/U202  ( .A0(\add_x_19_2/n162 ), .A1(\add_x_19_2/n166 ), 
        .B0(\add_x_19_2/n163 ), .Y(\add_x_19_2/n161 ) );
  XOR2X1TS \add_x_22_2/U72  ( .A(\add_x_22_2/n65 ), .B(\add_x_22_2/n64 ), .Y(
        \addr_calc/fir_read_calc/counter/N58 ) );
  NAND2X1TS \add_x_22_2/U81  ( .A(\add_x_22_2/n68 ), .B(n1690), .Y(
        \add_x_22_2/n65 ) );
  XNOR2X1TS \add_x_22_5/U47  ( .A(\add_x_22_5/n41 ), .B(n2047), .Y(
        \addr_calc/iir_write_calc/counter/N63 ) );
  NAND2X1TS \add_x_19_1/U102  ( .A(\add_x_19_1/n204 ), .B(\add_x_19_1/n98 ), 
        .Y(\add_x_19_1/n13 ) );
  XNOR2X1TS \add_x_22_1/U16  ( .A(\add_x_22_1/n16 ), .B(\add_x_22_1/n15 ), .Y(
        \addr_calc/fft_write_calc/counter/N69 ) );
  NOR2X1TS \add_x_19_1/U131  ( .A(\add_x_19_1/n135 ), .B(\add_x_19_1/n116 ), 
        .Y(\add_x_19_1/n114 ) );
  OAI21X1TS \add_x_19_1/U132  ( .A0(\add_x_19_1/n136 ), .A1(\add_x_19_1/n116 ), 
        .B0(\add_x_19_1/n117 ), .Y(\add_x_19_1/n115 ) );
  AOI21X1TS \add_x_19_1/U134  ( .A0(\add_x_19_1/n118 ), .A1(\add_x_19_1/n127 ), 
        .B0(\add_x_19_1/n119 ), .Y(\add_x_19_1/n117 ) );
  OAI21X1TS \add_x_19_1/U136  ( .A0(\add_x_19_1/n120 ), .A1(\add_x_19_1/n124 ), 
        .B0(\add_x_19_1/n121 ), .Y(\add_x_19_1/n119 ) );
  OAI21X1TS \add_x_19_1/U202  ( .A0(\add_x_19_1/n162 ), .A1(\add_x_19_1/n166 ), 
        .B0(\add_x_19_1/n163 ), .Y(\add_x_19_1/n161 ) );
  XNOR2X1TS \add_x_22_1/U126  ( .A(\add_x_22_1/n106 ), .B(n1158), .Y(
        \addr_calc/fft_write_calc/counter/N48 ) );
  NAND2X1TS \add_x_19_1/U217  ( .A(\add_x_19_1/n218 ), .B(\add_x_19_1/n171 ), 
        .Y(\add_x_19_1/n27 ) );
  TBUFX8TS \addr_calc/addr_tri3[15]  ( .A(\addr_calc/fir_read_addr[15] ), .OE(
        n2755), .Y(addr[15]) );
  TBUFX6TS \addr_calc/addr_tri[19]  ( .A(\addr_calc/fft_read_addr[19] ), .OE(
        n2738), .Y(addr[19]) );
  DFFHQX1TS \addr_calc/fir_read_calc/counter/count_reg[21]  ( .D(n1077), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[21] ) );
  TBUFX6TS \addr_calc/addr_tri5[15]  ( .A(\addr_calc/iir_read_addr[15] ), .OE(
        n2771), .Y(addr[15]) );
  TBUFX6TS \addr_calc/addr_tri4[28]  ( .A(\addr_calc/fir_write_addr[28] ), 
        .OE(n2759), .Y(addr[28]) );
  DFFHQX2TS \addr_calc/fft_write_calc/counter/count_reg[5]  ( .D(n1061), .CK(
        clk), .Q(\addr_calc/fft_write_calc/count[5] ) );
  TBUFX12TS \addr_calc/addr_tri3[25]  ( .A(\addr_calc/fir_read_addr[25] ), 
        .OE(n2752), .Y(addr[25]) );
  TBUFX4TS \addr_calc/addr_tri2[22]  ( .A(\addr_calc/fft_write_addr[22] ), 
        .OE(n2745), .Y(addr[22]) );
  TBUFX4TS \addr_calc/addr_tri5[13]  ( .A(\addr_calc/iir_read_addr[13] ), .OE(
        n2771), .Y(addr[13]) );
  TBUFX4TS \addr_calc/addr_tri3[13]  ( .A(\addr_calc/fir_read_addr[13] ), .OE(
        n2755), .Y(addr[13]) );
  TBUFX12TS \addr_calc/addr_tri3[28]  ( .A(\addr_calc/fir_read_addr[28] ), 
        .OE(n2751), .Y(addr[28]) );
  TBUFX16TS \addr_calc/addr_tri5[23]  ( .A(\addr_calc/iir_read_addr[23] ), 
        .OE(n2769), .Y(addr[23]) );
  TBUFX6TS \addr_calc/addr_tri[15]  ( .A(\addr_calc/fft_read_addr[15] ), .OE(
        n2739), .Y(addr[15]) );
  DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[11]  ( .D(n991), .CK(
        clk), .Q(\addr_calc/iir_write_calc/count[11] ) );
  TBUFX8TS \addr_calc/addr_tri2[19]  ( .A(\addr_calc/fft_write_addr[19] ), 
        .OE(n2746), .Y(addr[19]) );
  TBUFX16TS \addr_calc/addr_tri3[19]  ( .A(\addr_calc/fir_read_addr[19] ), 
        .OE(n2754), .Y(addr[19]) );
  TBUFX6TS \addr_calc/addr_tri4[25]  ( .A(\addr_calc/fir_write_addr[25] ), 
        .OE(n2760), .Y(addr[25]) );
  TBUFX12TS \addr_calc/addr_tri6[31]  ( .A(\addr_calc/iir_write_addr[31] ), 
        .OE(n2775), .Y(addr[31]) );
  TBUFX4TS \addr_calc/addr_tri3[17]  ( .A(\addr_calc/fir_read_addr[17] ), .OE(
        n2754), .Y(addr[17]) );
  TBUFX4TS \addr_calc/addr_tri3[20]  ( .A(\addr_calc/fir_read_addr[20] ), .OE(
        n2753), .Y(addr[20]) );
  TBUFX12TS \addr_calc/addr_tri2[25]  ( .A(\addr_calc/fft_write_addr[25] ), 
        .OE(n2744), .Y(addr[25]) );
  TBUFX12TS \addr_calc/addr_tri6[25]  ( .A(\addr_calc/iir_write_addr[25] ), 
        .OE(n2776), .Y(addr[25]) );
  TBUFX12TS \addr_calc/addr_tri6[28]  ( .A(\addr_calc/iir_write_addr[28] ), 
        .OE(n2775), .Y(addr[28]) );
  TBUFX8TS \addr_calc/addr_tri3[27]  ( .A(\addr_calc/fir_read_addr[27] ), .OE(
        n2752), .Y(addr[27]) );
  TBUFX12TS \addr_calc/addr_tri[27]  ( .A(\addr_calc/fft_read_addr[27] ), .OE(
        n2736), .Y(addr[27]) );
  TBUFX8TS \addr_calc/addr_tri6[27]  ( .A(\addr_calc/iir_write_addr[27] ), 
        .OE(n2776), .Y(addr[27]) );
  DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[9]  ( .D(n1089), .CK(
        clk), .Q(\addr_calc/fir_read_calc/count[9] ) );
  TBUFX12TS \addr_calc/addr_tri2[23]  ( .A(\addr_calc/fft_write_addr[23] ), 
        .OE(n2745), .Y(addr[23]) );
  TBUFX12TS \addr_calc/addr_tri2[31]  ( .A(\addr_calc/fft_write_addr[31] ), 
        .OE(n2743), .Y(addr[31]) );
  DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[6]  ( .D(n1028), .CK(
        clk), .Q(\addr_calc/fft_read_calc/count[6] ) );
  TBUFX16TS \addr_calc/addr_tri2[27]  ( .A(\addr_calc/fft_write_addr[27] ), 
        .OE(n2744), .Y(addr[27]) );
  TBUFX4TS \addr_calc/addr_tri5[29]  ( .A(\addr_calc/iir_read_addr[29] ), .OE(
        n2767), .Y(addr[29]) );
  INVX2TS U396 ( .A(n2795), .Y(n1720) );
  INVX4TS U397 ( .A(n2795), .Y(n1700) );
  INVX2TS U398 ( .A(n1720), .Y(n1727) );
  NAND2X8TS U399 ( .A(n1779), .B(n1780), .Y(
        \addr_calc/iir_write_calc/counter/N38 ) );
  XNOR2X2TS U400 ( .A(\add_x_19_3/n38 ), .B(n1538), .Y(
        \addr_calc/fir_write_addr[30] ) );
  OAI21X1TS U401 ( .A0(\add_x_19_4/n102 ), .A1(\add_x_19_4/n100 ), .B0(
        \add_x_19_4/n101 ), .Y(\add_x_19_4/n99 ) );
  XNOR2X2TS U402 ( .A(\DP_OP_158_296_6262/n841 ), .B(n1988), .Y(
        \DP_OP_158_296_6262/n202 ) );
  BUFX4TS U403 ( .A(n2660), .Y(n2655) );
  NOR2X2TS U404 ( .A(\add_x_19_0/n86 ), .B(\add_x_19_0/n89 ), .Y(
        \add_x_19_0/n84 ) );
  XOR2X4TS U405 ( .A(\add_x_19_2/n99 ), .B(n1137), .Y(
        \addr_calc/fir_read_addr[19] ) );
  AND2X6TS U406 ( .A(\add_x_19_2/n204 ), .B(\add_x_19_2/n98 ), .Y(n1137) );
  XOR2X4TS U407 ( .A(n1702), .B(n1971), .Y(\DP_OP_159_297_3515/n495 ) );
  NAND2X2TS U408 ( .A(\addr_calc/fft_read_calc/count[20] ), .B(n2440), .Y(
        \add_x_19_0/n90 ) );
  NOR2XLTS U409 ( .A(n1505), .B(n1510), .Y(n1138) );
  INVX1TS U410 ( .A(n1504), .Y(n1505) );
  AO22X4TS U411 ( .A0(n1761), .A1(\addr_calc/fir_write_calc/counter/N68 ), 
        .B0(n1894), .B1(n1259), .Y(n1105) );
  CLKINVX4TS U412 ( .A(n2803), .Y(n1757) );
  CLKINVX4TS U413 ( .A(n2803), .Y(n1758) );
  NOR2X4TS U414 ( .A(n1241), .B(n785), .Y(n2803) );
  INVX1TS U415 ( .A(\add_x_19_1/n92 ), .Y(\add_x_19_1/n91 ) );
  CLKINVX2TS U416 ( .A(\add_x_19_1/n69 ), .Y(\add_x_19_1/n68 ) );
  AOI21X2TS U417 ( .A0(\add_x_19_1/n112 ), .A1(\add_x_19_1/n103 ), .B0(
        \add_x_19_1/n104 ), .Y(\add_x_19_1/n102 ) );
  CLKXOR2X2TS U418 ( .A(\add_x_19_1/n68 ), .B(n1406), .Y(
        \addr_calc/fft_write_addr[24] ) );
  OAI21X1TS U419 ( .A0(\add_x_19_1/n60 ), .A1(\add_x_19_1/n58 ), .B0(
        \add_x_19_1/n59 ), .Y(\add_x_19_1/n57 ) );
  OAI2BB1X2TS U420 ( .A0N(n1552), .A1N(\add_x_19_1/n38 ), .B0(n1553), .Y(n1551) );
  OAI2BB1X2TS U421 ( .A0N(n2052), .A1N(n2655), .B0(n1608), .Y(n1028) );
  INVX2TS U422 ( .A(n1700), .Y(n1694) );
  BUFX3TS U423 ( .A(\add_x_19_0/n113 ), .Y(n1139) );
  XOR2XLTS U424 ( .A(\add_x_19_0/n91 ), .B(n1393), .Y(
        \addr_calc/fft_read_addr[20] ) );
  MXI2X4TS U425 ( .A(n2798), .B(\addr_calc/fft_write_calc/counter/N43 ), .S0(
        n2662), .Y(n1066) );
  XOR2X4TS U426 ( .A(n1731), .B(\add_x_22_1/n30 ), .Y(
        \DP_OP_158_296_6262/n580 ) );
  XOR2X1TS U427 ( .A(\add_x_19_2/n60 ), .B(n1325), .Y(
        \addr_calc/fir_read_addr[26] ) );
  OAI2BB1X2TS U428 ( .A0N(n1229), .A1N(\add_x_19_2/n60 ), .B0(n1230), .Y(n1228) );
  XOR2XLTS U429 ( .A(\add_x_19_2/n156 ), .B(\add_x_19_2/n24 ), .Y(
        \addr_calc/fir_read_addr[8] ) );
  XOR2X4TS U430 ( .A(\add_x_19_3/n35 ), .B(n1140), .Y(
        \addr_calc/fir_write_addr[31] ) );
  AND2X6TS U431 ( .A(n2630), .B(\add_x_19_3/n34 ), .Y(n1140) );
  CLKINVX4TS U432 ( .A(n1701), .Y(n1751) );
  NAND2X1TS U433 ( .A(n1826), .B(\addr_calc/fir_read_calc/counter/N47 ), .Y(
        n1141) );
  NAND2XLTS U434 ( .A(n1663), .B(n1906), .Y(n1142) );
  NAND2X1TS U435 ( .A(n1141), .B(n1142), .Y(n1094) );
  INVX3TS U436 ( .A(n2809), .Y(n1742) );
  AOI21X1TS U437 ( .A0(\add_x_19_5/n92 ), .A1(\add_x_19_5/n84 ), .B0(
        \add_x_19_5/n85 ), .Y(\add_x_19_5/n83 ) );
  NOR2X2TS U438 ( .A(\DP_OP_159_297_3515/n1026 ), .B(
        \DP_OP_159_297_3515/n1014 ), .Y(\DP_OP_159_297_3515/n1011 ) );
  AOI21X2TS U439 ( .A0(\add_x_19_4/n127 ), .A1(n1549), .B0(\add_x_19_4/n119 ), 
        .Y(\add_x_19_4/n117 ) );
  CLKINVX3TS U440 ( .A(n1897), .Y(n1540) );
  NAND4BXLTS U441 ( .AN(\add_x_22_2/n103 ), .B(\add_x_22_2/n111 ), .C(
        \addr_calc/fir_read_calc/count[7] ), .D(n2001), .Y(\add_x_22_2/n94 )
         );
  XNOR2X4TS U442 ( .A(n1596), .B(n1597), .Y(\addr_calc/fir_read_addr[23] ) );
  OAI21X1TS U443 ( .A0(\add_x_19_1/n83 ), .A1(\add_x_19_1/n81 ), .B0(
        \add_x_19_1/n82 ), .Y(\add_x_19_1/n80 ) );
  NOR4BBX1TS U444 ( .AN(n1899), .BN(n1143), .C(n1480), .D(n2001), .Y(n877) );
  INVX20TS U445 ( .A(n1997), .Y(n1143) );
  AOI2BB1X2TS U446 ( .A0N(\add_x_19_2/n60 ), .A1N(n1227), .B0(n1228), .Y(
        \addr_calc/fir_read_addr[27] ) );
  AOI21X1TS U447 ( .A0(\add_x_19_1/n69 ), .A1(\add_x_19_1/n61 ), .B0(
        \add_x_19_1/n62 ), .Y(\add_x_19_1/n60 ) );
  BUFX2TS U448 ( .A(\DP_OP_158_296_6262/n1999 ), .Y(n1144) );
  NAND2X6TS U449 ( .A(\DP_OP_158_296_6262/n1986 ), .B(
        \DP_OP_158_296_6262/n1931 ), .Y(n2589) );
  CLKINVX2TS U450 ( .A(n1720), .Y(n1145) );
  CLKINVX1TS U451 ( .A(n1700), .Y(n1726) );
  NOR2X2TS U452 ( .A(n1892), .B(n2450), .Y(\add_x_19_3/n86 ) );
  INVX3TS U453 ( .A(n1891), .Y(n1892) );
  AND2X6TS U454 ( .A(n1789), .B(\DP_OP_159_297_3515/n963 ), .Y(n1698) );
  CLKINVX4TS U455 ( .A(n2047), .Y(n2048) );
  NOR2X4TS U456 ( .A(\DP_OP_159_297_3515/n971 ), .B(\DP_OP_159_297_3515/n959 ), 
        .Y(\DP_OP_159_297_3515/n956 ) );
  XOR2X4TS U457 ( .A(\DP_OP_158_296_6262/n1950 ), .B(\DP_OP_159_297_3515/n871 ), .Y(n1659) );
  CLKINVX2TS U458 ( .A(n1503), .Y(\DP_OP_159_297_3515/n871 ) );
  XNOR2X2TS U459 ( .A(n2621), .B(\addr_calc/iir_read_calc/count[10] ), .Y(
        \DP_OP_159_297_3515/n289 ) );
  NOR2X2TS U460 ( .A(\DP_OP_159_297_3515/n1052 ), .B(
        \DP_OP_159_297_3515/n1041 ), .Y(\DP_OP_159_297_3515/n1040 ) );
  NAND2X2TS U461 ( .A(\DP_OP_158_296_6262/n320 ), .B(\DP_OP_158_296_6262/n347 ), .Y(\DP_OP_158_296_6262/n318 ) );
  NOR2X4TS U462 ( .A(\DP_OP_158_296_6262/n1171 ), .B(
        \DP_OP_158_296_6262/n1160 ), .Y(\DP_OP_158_296_6262/n1158 ) );
  CLKINVX3TS U463 ( .A(n1782), .Y(n1789) );
  CLKINVX2TS U464 ( .A(\add_x_19_4/n92 ), .Y(\add_x_19_4/n91 ) );
  BUFX6TS U465 ( .A(n2670), .Y(n2668) );
  XOR2X1TS U466 ( .A(\add_x_19_2/n91 ), .B(n1404), .Y(
        \addr_calc/fir_read_addr[20] ) );
  XNOR2XLTS U467 ( .A(n1635), .B(\addr_calc/fft_read_calc/count[17] ), .Y(
        n1634) );
  INVXLTS U468 ( .A(\add_x_19_0/n105 ), .Y(\add_x_19_0/n206 ) );
  XNOR2X1TS U469 ( .A(n2614), .B(n1847), .Y(\DP_OP_159_297_3515/n5 ) );
  XOR2X4TS U470 ( .A(\DP_OP_159_297_3515/n934 ), .B(n1146), .Y(n1738) );
  INVX20TS U471 ( .A(\DP_OP_158_296_6262/n1869 ), .Y(n1146) );
  XNOR2X2TS U472 ( .A(n1756), .B(n2023), .Y(\DP_OP_158_296_6262/n724 ) );
  AOI21X1TS U473 ( .A0(\add_x_19_1/n177 ), .A1(\add_x_19_1/n168 ), .B0(n1157), 
        .Y(\add_x_19_1/n167 ) );
  NOR2X2TS U474 ( .A(n2410), .B(n1999), .Y(\add_x_19_3/n131 ) );
  INVX4TS U475 ( .A(n1998), .Y(n1999) );
  OAI21X2TS U476 ( .A0(\add_x_19_3/n68 ), .A1(\add_x_19_3/n66 ), .B0(
        \add_x_19_3/n67 ), .Y(\add_x_19_3/n65 ) );
  INVX1TS U477 ( .A(\add_x_19_0/n72 ), .Y(\add_x_19_0/n70 ) );
  CLKINVX8TS U478 ( .A(n2589), .Y(n1793) );
  XNOR2X4TS U479 ( .A(n1356), .B(n1357), .Y(\addr_calc/iir_read_addr[31] ) );
  NAND2XLTS U480 ( .A(\DP_OP_158_296_6262/n1959 ), .B(
        \DP_OP_158_296_6262/n1945 ), .Y(\DP_OP_158_296_6262/n1944 ) );
  OAI21XLTS U481 ( .A0(n2793), .A1(n2057), .B0(fft_enable), .Y(n1394) );
  XNOR2X1TS U482 ( .A(\add_x_19_5/n65 ), .B(\add_x_19_5/n7 ), .Y(
        \addr_calc/iir_write_addr[25] ) );
  NOR2BX2TS U483 ( .AN(n1632), .B(\add_x_19_4/n131 ), .Y(\add_x_19_4/n126 ) );
  INVX2TS U484 ( .A(\add_x_19_4/n73 ), .Y(\add_x_19_4/n71 ) );
  OAI21X2TS U485 ( .A0(\add_x_19_4/n132 ), .A1(\add_x_19_4/n128 ), .B0(
        \add_x_19_4/n129 ), .Y(\add_x_19_4/n127 ) );
  XNOR2X1TS U486 ( .A(n1776), .B(n2017), .Y(\DP_OP_158_296_6262/n621 ) );
  NAND2X2TS U487 ( .A(n1677), .B(n1462), .Y(n1147) );
  XOR2X4TS U488 ( .A(n1730), .B(n1949), .Y(\DP_OP_158_296_6262/n1027 ) );
  CLKINVX1TS U489 ( .A(n1509), .Y(n1511) );
  INVX1TS U490 ( .A(n1509), .Y(n1510) );
  CLKINVX2TS U491 ( .A(\DP_OP_158_296_6262/n1958 ), .Y(
        \DP_OP_158_296_6262/n1959 ) );
  XOR2X4TS U492 ( .A(n1777), .B(n1841), .Y(\DP_OP_158_296_6262/n39 ) );
  OAI21X2TS U493 ( .A0(\add_x_19_3/n68 ), .A1(\add_x_19_3/n51 ), .B0(
        \add_x_19_3/n52 ), .Y(\add_x_19_3/n50 ) );
  AOI21X2TS U494 ( .A0(\add_x_19_5/n137 ), .A1(\add_x_19_5/n150 ), .B0(
        \add_x_19_5/n138 ), .Y(\add_x_19_5/n136 ) );
  NAND2X2TS U495 ( .A(\DP_OP_158_296_6262/n1973 ), .B(n1591), .Y(
        \DP_OP_158_296_6262/n1958 ) );
  XOR2X2TS U496 ( .A(\add_x_19_0/n57 ), .B(n1465), .Y(
        \addr_calc/fft_read_addr[27] ) );
  XNOR2X2TS U497 ( .A(n1658), .B(\addr_calc/fft_read_calc/count[15] ), .Y(
        \DP_OP_158_296_6262/n1136 ) );
  NOR2X6TS U498 ( .A(\DP_OP_158_296_6262/n998 ), .B(\DP_OP_158_296_6262/n1013 ), .Y(\DP_OP_158_296_6262/n996 ) );
  MXI2X4TS U499 ( .A(\DP_OP_159_297_3515/n880 ), .B(\DP_OP_159_297_3515/n1066 ), .S0(\DP_OP_159_297_3515/n1075 ), .Y(\DP_OP_159_297_3515/n1064 ) );
  XNOR2X4TS U500 ( .A(n2620), .B(n1942), .Y(\DP_OP_159_297_3515/n705 ) );
  NAND2X4TS U501 ( .A(n1734), .B(n1735), .Y(n2620) );
  NOR2X4TS U502 ( .A(n1516), .B(n1518), .Y(\DP_OP_158_296_6262/n1878 ) );
  CLKINVX2TS U503 ( .A(n1517), .Y(n1518) );
  NOR2X2TS U504 ( .A(\DP_OP_158_296_6262/n702 ), .B(\DP_OP_158_296_6262/n689 ), 
        .Y(\DP_OP_158_296_6262/n687 ) );
  INVX1TS U505 ( .A(n1526), .Y(n1527) );
  XNOR2X2TS U506 ( .A(n1651), .B(n1666), .Y(\DP_OP_158_296_6262/n1216 ) );
  NOR2X4TS U507 ( .A(n2424), .B(\addr_calc/iir_read_calc/count[14] ), .Y(
        \add_x_19_4/n123 ) );
  NOR2X2TS U508 ( .A(n1911), .B(n2404), .Y(\add_x_19_4/n139 ) );
  XOR2X4TS U509 ( .A(n1147), .B(n1484), .Y(n1655) );
  NOR2X4TS U510 ( .A(n1503), .B(n1457), .Y(\DP_OP_158_296_6262/n1945 ) );
  OAI31X1TS U511 ( .A0(\add_x_19_3/n128 ), .A1(n1300), .A2(n1301), .B0(n1302), 
        .Y(\addr_calc/fir_write_addr[13] ) );
  NAND2X2TS U512 ( .A(\add_x_19_2/n168 ), .B(\add_x_19_2/n160 ), .Y(
        \add_x_19_2/n158 ) );
  XNOR2X4TS U513 ( .A(\add_x_19_4/n50 ), .B(\add_x_19_4/n4 ), .Y(
        \addr_calc/iir_read_addr[28] ) );
  XNOR2X4TS U514 ( .A(\add_x_19_4/n65 ), .B(\add_x_19_4/n7 ), .Y(
        \addr_calc/iir_read_addr[25] ) );
  NAND4XLTS U515 ( .A(n876), .B(n877), .C(n878), .D(n879), .Y(n2799) );
  NOR4X1TS U516 ( .A(n1838), .B(n2004), .C(n1842), .D(n1871), .Y(n879) );
  INVX3TS U517 ( .A(n1870), .Y(n1871) );
  NOR2X2TS U518 ( .A(n1683), .B(n2420), .Y(\add_x_19_5/n162 ) );
  INVX2TS U519 ( .A(n1938), .Y(n1683) );
  OAI21X1TS U520 ( .A0(\add_x_19_0/n60 ), .A1(\add_x_19_0/n58 ), .B0(
        \add_x_19_0/n59 ), .Y(\add_x_19_0/n57 ) );
  NOR2X4TS U521 ( .A(\DP_OP_158_296_6262/n515 ), .B(\DP_OP_158_296_6262/n534 ), 
        .Y(\DP_OP_158_296_6262/n513 ) );
  NAND2X2TS U522 ( .A(\addr_calc/fft_write_calc/count[5] ), .B(n2484), .Y(
        \add_x_19_1/n171 ) );
  XOR2XLTS U523 ( .A(\add_x_19_1/n156 ), .B(n1405), .Y(
        \addr_calc/fft_write_addr[8] ) );
  XNOR2XLTS U524 ( .A(n1447), .B(\add_x_19_1/n112 ), .Y(
        \addr_calc/fft_write_addr[16] ) );
  XNOR2XLTS U525 ( .A(n1446), .B(\add_x_19_1/n146 ), .Y(
        \addr_calc/fft_write_addr[10] ) );
  NOR2X2TS U526 ( .A(n1670), .B(n2489), .Y(\add_x_19_3/n97 ) );
  CLKINVX6TS U527 ( .A(n1889), .Y(n1670) );
  NOR2X2TS U528 ( .A(n1686), .B(n2483), .Y(\add_x_19_5/n170 ) );
  XNOR2X2TS U529 ( .A(\add_x_19_3/n80 ), .B(\add_x_19_3/n9 ), .Y(
        \addr_calc/fir_write_addr[23] ) );
  NAND2XLTS U530 ( .A(\add_x_22_3/n68 ), .B(
        \addr_calc/fir_write_calc/count[14] ), .Y(\add_x_22_3/n65 ) );
  OAI21X1TS U531 ( .A0(\add_x_19_3/n113 ), .A1(\add_x_19_3/n70 ), .B0(
        \add_x_19_3/n71 ), .Y(\add_x_19_3/n69 ) );
  NAND4BXLTS U532 ( .AN(\add_x_22_3/n69 ), .B(n2003), .C(n1883), .D(
        \add_x_22_3/n77 ), .Y(n1273) );
  OR2X6TS U533 ( .A(n2003), .B(n2426), .Y(n1545) );
  INVX3TS U534 ( .A(\addr_calc/fir_write_calc/count[14] ), .Y(n2002) );
  INVX1TS U535 ( .A(n1512), .Y(n1457) );
  INVX3TS U536 ( .A(\addr_calc/fir_write_calc/count[19] ), .Y(n1889) );
  CLKINVX2TS U537 ( .A(\addr_calc/fft_read_calc/count[20] ), .Y(
        \add_x_22_0/n40 ) );
  NOR2BX2TS U538 ( .AN(n2439), .B(\addr_calc/fft_read_calc/count[20] ), .Y(
        \add_x_19_0/n89 ) );
  NOR2X4TS U539 ( .A(n1905), .B(n2420), .Y(\add_x_19_4/n162 ) );
  CLKINVX4TS U540 ( .A(\addr_calc/fft_write_calc/count[5] ), .Y(n1158) );
  NOR2X2TS U541 ( .A(n1728), .B(n2364), .Y(\DP_OP_158_296_6262/n1978 ) );
  NOR2X2TS U542 ( .A(n1728), .B(\DP_OP_158_296_6262/n1972 ), .Y(
        \DP_OP_158_296_6262/n1971 ) );
  NOR2X2TS U543 ( .A(n1728), .B(\DP_OP_158_296_6262/n1937 ), .Y(
        \DP_OP_158_296_6262/n1936 ) );
  CLKINVX2TS U544 ( .A(n1511), .Y(\DP_OP_159_297_3515/n875 ) );
  INVX1TS U545 ( .A(n2482), .Y(n2484) );
  INVX2TS U546 ( .A(n1742), .Y(n1674) );
  INVX3TS U547 ( .A(n1899), .Y(n1900) );
  CLKINVX1TS U548 ( .A(n1819), .Y(n1148) );
  XOR2X4TS U549 ( .A(n1736), .B(n1678), .Y(n1149) );
  XOR2XLTS U550 ( .A(\add_x_19_1/n91 ), .B(n1441), .Y(
        \addr_calc/fft_write_addr[20] ) );
  XOR2X4TS U551 ( .A(\DP_OP_158_296_6262/n833 ), .B(\add_x_22_1/n15 ), .Y(
        \DP_OP_158_296_6262/n534 ) );
  XNOR2X1TS U552 ( .A(\add_x_19_1/n60 ), .B(n1150), .Y(
        \addr_calc/fft_write_addr[26] ) );
  INVX20TS U553 ( .A(n1321), .Y(n1150) );
  CLKINVX3TS U554 ( .A(n1700), .Y(n1721) );
  AO22X4TS U555 ( .A0(n1823), .A1(\addr_calc/fir_read_calc/counter/N59 ), .B0(
        n1743), .B1(\addr_calc/fir_read_calc/count[16] ), .Y(n1082) );
  AO22X4TS U556 ( .A0(n1823), .A1(\addr_calc/fir_read_calc/counter/N61 ), .B0(
        n1743), .B1(\addr_calc/fir_read_calc/count[18] ), .Y(n1080) );
  NAND2BX2TS U557 ( .AN(n2047), .B(n2441), .Y(\add_x_19_5/n90 ) );
  NAND2XLTS U558 ( .A(n1489), .B(n1506), .Y(\DP_OP_159_297_3515/n1041 ) );
  XNOR2X2TS U559 ( .A(n2619), .B(n1785), .Y(\DP_OP_159_297_3515/n269 ) );
  CLKINVX1TS U560 ( .A(n1504), .Y(n1506) );
  INVXLTS U561 ( .A(\add_x_19_0/n134 ), .Y(\add_x_19_0/n133 ) );
  BUFX8TS U562 ( .A(n2807), .Y(n1151) );
  OAI2BB1XLTS U563 ( .A0N(n1822), .A1N(\addr_calc/fir_read_calc/counter/N73 ), 
        .B0(n1645), .Y(n1068) );
  BUFX4TS U564 ( .A(n2803), .Y(n1152) );
  NAND2BXLTS U565 ( .AN(n1189), .B(n1822), .Y(n1188) );
  AO22X2TS U566 ( .A0(n1821), .A1(\addr_calc/fir_read_calc/counter/N50 ), .B0(
        n1743), .B1(n1480), .Y(n1091) );
  NAND2BXLTS U567 ( .AN(n1203), .B(n1148), .Y(n1202) );
  AO22X2TS U568 ( .A0(n1826), .A1(\addr_calc/fir_read_calc/counter/N44 ), .B0(
        n1672), .B1(n1910), .Y(n1097) );
  NAND2BX1TS U569 ( .AN(n1168), .B(n1826), .Y(n1167) );
  AO22X2TS U570 ( .A0(n1825), .A1(\addr_calc/fir_read_calc/counter/N48 ), .B0(
        n1672), .B1(n1904), .Y(n1093) );
  NAND2BXLTS U571 ( .AN(n1185), .B(n1825), .Y(n1184) );
  BUFX4TS U572 ( .A(n2660), .Y(n2656) );
  CLKINVX1TS U573 ( .A(n1512), .Y(n1513) );
  CLKINVX4TS U574 ( .A(n1474), .Y(n1475) );
  INVX3TS U575 ( .A(n1701), .Y(n1754) );
  CLKINVX3TS U576 ( .A(n1746), .Y(n1747) );
  CLKINVX3TS U577 ( .A(n1746), .Y(n1460) );
  OAI2BB1X1TS U578 ( .A0N(n1873), .A1N(n1747), .B0(n1202), .Y(n1071) );
  INVX4TS U579 ( .A(n1758), .Y(n1762) );
  CLKINVX4TS U580 ( .A(n1474), .Y(n1477) );
  CLKINVX2TS U581 ( .A(n2795), .Y(n1719) );
  CLKINVX3TS U582 ( .A(n1700), .Y(n1722) );
  CLKINVX4TS U583 ( .A(n2807), .Y(n1820) );
  XNOR2X4TS U584 ( .A(n1652), .B(n1665), .Y(\DP_OP_158_296_6262/n1042 ) );
  NOR2X4TS U585 ( .A(n1523), .B(n1531), .Y(\DP_OP_158_296_6262/n1906 ) );
  CLKINVX8TS U586 ( .A(n1741), .Y(n1746) );
  NAND2X4TS U587 ( .A(\DP_OP_158_296_6262/n606 ), .B(\DP_OP_158_296_6262/n578 ), .Y(\DP_OP_158_296_6262/n576 ) );
  INVX1TS U588 ( .A(n1158), .Y(n1479) );
  OAI21XLTS U589 ( .A0(\add_x_19_1/n170 ), .A1(\add_x_19_1/n176 ), .B0(
        \add_x_19_1/n171 ), .Y(n1157) );
  OAI21X2TS U590 ( .A0(\add_x_19_1/n170 ), .A1(\add_x_19_1/n176 ), .B0(
        \add_x_19_1/n171 ), .Y(\add_x_19_1/n169 ) );
  AOI21X4TS U591 ( .A0(\add_x_19_1/n157 ), .A1(\add_x_19_1/n114 ), .B0(
        \add_x_19_1/n115 ), .Y(\add_x_19_1/n113 ) );
  OAI21X2TS U592 ( .A0(\add_x_19_1/n113 ), .A1(\add_x_19_1/n93 ), .B0(
        \add_x_19_1/n94 ), .Y(\add_x_19_1/n92 ) );
  OAI21X2TS U593 ( .A0(\add_x_19_1/n44 ), .A1(\add_x_19_1/n113 ), .B0(
        \add_x_19_1/n45 ), .Y(\add_x_19_1/n43 ) );
  INVX2TS U594 ( .A(\add_x_19_1/n113 ), .Y(\add_x_19_1/n112 ) );
  OAI21X2TS U595 ( .A0(\add_x_19_1/n113 ), .A1(\add_x_19_1/n70 ), .B0(
        \add_x_19_1/n71 ), .Y(\add_x_19_1/n69 ) );
  AOI21X2TS U596 ( .A0(\add_x_19_1/n92 ), .A1(\add_x_19_1/n84 ), .B0(
        \add_x_19_1/n85 ), .Y(\add_x_19_1/n83 ) );
  XNOR2X1TS U597 ( .A(\add_x_19_1/n83 ), .B(n1154), .Y(
        \addr_calc/fft_write_addr[22] ) );
  NAND2BX1TS U598 ( .AN(\add_x_19_1/n81 ), .B(\add_x_19_1/n82 ), .Y(n1153) );
  INVX2TS U599 ( .A(n1153), .Y(n1154) );
  NAND2X2TS U600 ( .A(\DP_OP_158_296_6262/n2010 ), .B(n1144), .Y(
        \DP_OP_158_296_6262/n1998 ) );
  INVX2TS U601 ( .A(n1485), .Y(n1155) );
  NOR2X4TS U602 ( .A(\addr_calc/iir_read_calc/count[15] ), .B(n2475), .Y(
        \add_x_19_4/n120 ) );
  INVXLTS U603 ( .A(\add_x_19_1/n170 ), .Y(\add_x_19_1/n218 ) );
  XNOR2X1TS U604 ( .A(\add_x_19_4/n83 ), .B(n1156), .Y(
        \addr_calc/iir_read_addr[22] ) );
  INVX20TS U605 ( .A(n1433), .Y(n1156) );
  INVXLTS U606 ( .A(n1526), .Y(n2363) );
  XOR2X2TS U607 ( .A(n2595), .B(\addr_calc/fft_read_calc/count[5] ), .Y(n1602)
         );
  XNOR2X4TS U608 ( .A(n2607), .B(n1954), .Y(\DP_OP_159_297_3515/n638 ) );
  OR3X2TS U609 ( .A(\data_cntl/N191 ), .B(n2785), .C(n1860), .Y(n1737) );
  NOR2X4TS U610 ( .A(\DP_OP_159_297_3515/n1 ), .B(\DP_OP_159_297_3515/n160 ), 
        .Y(n1781) );
  XOR2X4TS U611 ( .A(n2625), .B(\addr_calc/iir_write_calc/count[30] ), .Y(
        n1564) );
  XOR2X4TS U612 ( .A(\DP_OP_159_297_3515/n1128 ), .B(
        \addr_calc/iir_write_calc/count[18] ), .Y(\DP_OP_159_297_3515/n625 )
         );
  NOR2X4TS U613 ( .A(n1520), .B(n1482), .Y(\DP_OP_158_296_6262/n1933 ) );
  BUFX6TS U614 ( .A(n2797), .Y(n2670) );
  XNOR2X2TS U615 ( .A(\add_x_19_5/n50 ), .B(\add_x_19_5/n4 ), .Y(
        \addr_calc/iir_write_addr[28] ) );
  NAND2BX1TS U616 ( .AN(n1158), .B(n1939), .Y(\add_x_22_1/n103 ) );
  AOI21X4TS U617 ( .A0(\add_x_19_1/n169 ), .A1(\add_x_19_1/n160 ), .B0(
        \add_x_19_1/n161 ), .Y(\add_x_19_1/n159 ) );
  OAI21X4TS U618 ( .A0(\add_x_19_1/n178 ), .A1(\add_x_19_1/n158 ), .B0(
        \add_x_19_1/n159 ), .Y(\add_x_19_1/n157 ) );
  INVX2TS U619 ( .A(\add_x_19_1/n157 ), .Y(\add_x_19_1/n156 ) );
  NAND2X2TS U620 ( .A(\add_x_19_1/n168 ), .B(\add_x_19_1/n160 ), .Y(
        \add_x_19_1/n158 ) );
  XNOR2X4TS U621 ( .A(n1161), .B(n1912), .Y(n1159) );
  NOR2BX4TS U622 ( .AN(\add_x_22_1/n16 ), .B(n1162), .Y(n1161) );
  INVX12TS U623 ( .A(n2574), .Y(n1162) );
  NAND2X1TS U624 ( .A(n2669), .B(\addr_calc/fft_write_calc/count[27] ), .Y(
        n1160) );
  OAI2BB1X2TS U625 ( .A0N(n1694), .A1N(n1159), .B0(n1160), .Y(n1039) );
  XNOR2X4TS U626 ( .A(\add_x_22_1/n23 ), .B(n1165), .Y(n1164) );
  INVX12TS U627 ( .A(n2010), .Y(n1165) );
  NAND2BX1TS U628 ( .AN(n1164), .B(n1721), .Y(n1163) );
  OAI2BB1X1TS U629 ( .A0N(n2668), .A1N(\addr_calc/fft_write_calc/count[24] ), 
        .B0(n1163), .Y(n1042) );
  NAND2X1TS U630 ( .A(n1723), .B(\addr_calc/fft_write_calc/counter/N69 ), .Y(
        n1166) );
  OAI2BB1X1TS U631 ( .A0N(n2574), .A1N(n2668), .B0(n1166), .Y(n1040) );
  XNOR2X4TS U632 ( .A(n1169), .B(n1875), .Y(n1168) );
  NAND2BX4TS U633 ( .AN(n1170), .B(\add_x_22_2/n23 ), .Y(n1169) );
  INVX12TS U634 ( .A(\addr_calc/fir_read_calc/count[24] ), .Y(n1170) );
  OAI2BB1X1TS U635 ( .A0N(\addr_calc/fir_read_calc/count[25] ), .A1N(n1460), 
        .B0(n1167), .Y(n1073) );
  XNOR2X4TS U636 ( .A(\add_x_22_3/n16 ), .B(n1173), .Y(n1172) );
  INVX12TS U637 ( .A(\add_x_22_3/n15 ), .Y(n1173) );
  NAND2BX1TS U638 ( .AN(n1172), .B(n1764), .Y(n1171) );
  OAI2BB1X1TS U639 ( .A0N(n2581), .A1N(n1259), .B0(n1171), .Y(n1104) );
  CLKINVX1TS U640 ( .A(\add_x_19_1/n97 ), .Y(\add_x_19_1/n204 ) );
  OAI21X1TS U641 ( .A0(\add_x_19_1/n102 ), .A1(\add_x_19_1/n100 ), .B0(
        \add_x_19_1/n101 ), .Y(\add_x_19_1/n99 ) );
  XNOR2X2TS U642 ( .A(\add_x_19_1/n99 ), .B(\add_x_19_1/n13 ), .Y(
        \addr_calc/fft_write_addr[19] ) );
  OAI2BB1X4TS U643 ( .A0N(\add_x_19_3/n59 ), .A1N(n1178), .B0(n1179), .Y(n1177) );
  OAI2BB1X4TS U644 ( .A0N(\add_x_19_3/n58 ), .A1N(\add_x_19_3/n59 ), .B0(n1180), .Y(n1179) );
  INVX12TS U645 ( .A(n1178), .Y(n1180) );
  NOR2BX4TS U646 ( .AN(\add_x_19_3/n59 ), .B(n1178), .Y(n1176) );
  NAND2BX4TS U647 ( .AN(\add_x_19_3/n58 ), .B(n1178), .Y(n1174) );
  NOR2BX4TS U648 ( .AN(\add_x_19_3/n56 ), .B(\add_x_19_3/n55 ), .Y(n1178) );
  AOI2BB1X2TS U649 ( .A0N(\add_x_19_3/n60 ), .A1N(n1174), .B0(n1175), .Y(
        \addr_calc/fir_write_addr[27] ) );
  OAI2BB1X4TS U650 ( .A0N(n1176), .A1N(\add_x_19_3/n60 ), .B0(n1177), .Y(n1175) );
  XNOR2X4TS U651 ( .A(\add_x_22_5/n50 ), .B(n1183), .Y(n1182) );
  INVX12TS U652 ( .A(\add_x_22_5/n49 ), .Y(n1183) );
  NAND2BX1TS U653 ( .AN(n1182), .B(n1767), .Y(n1181) );
  OAI2BB1X2TS U654 ( .A0N(n2571), .A1N(n2676), .B0(n1181), .Y(n984) );
  AO22X4TS U655 ( .A0(n1768), .A1(\addr_calc/iir_write_calc/counter/N63 ), 
        .B0(n2676), .B1(\addr_calc/iir_write_calc/count[20] ), .Y(n982) );
  XNOR2X4TS U656 ( .A(n1186), .B(\add_x_22_2/n114 ), .Y(n1185) );
  NAND2BX4TS U657 ( .AN(n1187), .B(\add_x_22_2/n118 ), .Y(n1186) );
  INVX12TS U658 ( .A(n2004), .Y(n1187) );
  OAI2BB1X1TS U659 ( .A0N(n1908), .A1N(n1460), .B0(n1184), .Y(n1095) );
  AO22X2TS U660 ( .A0(n1148), .A1(\addr_calc/fir_read_calc/counter/N58 ), .B0(
        n1663), .B1(n1890), .Y(n1083) );
  XNOR2X4TS U661 ( .A(\add_x_22_2/n1 ), .B(n2549), .Y(n1189) );
  OAI2BB1X1TS U662 ( .A0N(n2549), .A1N(n1747), .B0(n1188), .Y(n1132) );
  INVX12TS U663 ( .A(\addr_calc/fir_write_calc/counter/N58 ), .Y(n1191) );
  NAND2BX1TS U664 ( .AN(n1191), .B(n1764), .Y(n1190) );
  OAI2BB1X2TS U665 ( .A0N(\addr_calc/fir_write_calc/count[15] ), .A1N(n1260), 
        .B0(n1190), .Y(n1115) );
  NOR2X2TS U666 ( .A(\add_x_19_2/n162 ), .B(\add_x_19_2/n165 ), .Y(
        \add_x_19_2/n160 ) );
  OAI21X1TS U667 ( .A0(\add_x_19_2/n136 ), .A1(\add_x_19_2/n116 ), .B0(
        \add_x_19_2/n117 ), .Y(\add_x_19_2/n115 ) );
  AOI21X4TS U668 ( .A0(\add_x_19_2/n157 ), .A1(\add_x_19_2/n114 ), .B0(
        \add_x_19_2/n115 ), .Y(\add_x_19_2/n113 ) );
  INVX1TS U669 ( .A(\add_x_19_2/n73 ), .Y(\add_x_19_2/n71 ) );
  INVX1TS U670 ( .A(\add_x_19_2/n72 ), .Y(\add_x_19_2/n70 ) );
  OAI21X2TS U671 ( .A0(\add_x_19_2/n113 ), .A1(\add_x_19_2/n70 ), .B0(
        \add_x_19_2/n71 ), .Y(\add_x_19_2/n69 ) );
  CLKINVX1TS U672 ( .A(\add_x_19_2/n63 ), .Y(\add_x_19_2/n198 ) );
  XNOR2X2TS U673 ( .A(\add_x_19_2/n65 ), .B(\add_x_19_2/n7 ), .Y(
        \addr_calc/fir_read_addr[25] ) );
  INVX1TS U674 ( .A(\add_x_19_2/n48 ), .Y(\add_x_19_2/n195 ) );
  XNOR2X2TS U675 ( .A(\add_x_19_2/n50 ), .B(\add_x_19_2/n4 ), .Y(
        \addr_calc/fir_read_addr[28] ) );
  AOI21X4TS U676 ( .A0(\addr_calc/iir_read_calc/counter/N38 ), .A1(data_to_iir), .B0(n1860), .Y(n2654) );
  AOI21X4TS U677 ( .A0(\addr_calc/iir_read_calc/counter/N38 ), .A1(data_to_iir), .B0(n1860), .Y(n1192) );
  BUFX4TS U678 ( .A(n1192), .Y(n1193) );
  BUFX6TS U679 ( .A(n1192), .Y(n2648) );
  BUFX6TS U680 ( .A(n1192), .Y(n2650) );
  BUFX4TS U681 ( .A(n1192), .Y(n2651) );
  AO22X2TS U682 ( .A0(n1714), .A1(\addr_calc/iir_read_calc/counter/N49 ), .B0(
        n1193), .B1(n2018), .Y(n965) );
  AO22X2TS U683 ( .A0(n1707), .A1(\addr_calc/iir_read_calc/counter/N47 ), .B0(
        n1193), .B1(n1903), .Y(n967) );
  AO22X4TS U684 ( .A0(n1710), .A1(\addr_calc/iir_read_calc/counter/N46 ), .B0(
        n1193), .B1(\addr_calc/iir_read_calc/count[3] ), .Y(n968) );
  AO22X4TS U685 ( .A0(n1712), .A1(\addr_calc/iir_read_calc/counter/N48 ), .B0(
        n1193), .B1(n2553), .Y(n966) );
  INVX12TS U686 ( .A(\addr_calc/iir_read_calc/counter/N64 ), .Y(n1195) );
  NAND2BX2TS U687 ( .AN(n1195), .B(n1712), .Y(n1194) );
  OAI2BB1X2TS U688 ( .A0N(\addr_calc/iir_read_calc/count[21] ), .A1N(n2652), 
        .B0(n1194), .Y(n950) );
  NAND2BX1TS U689 ( .AN(n2786), .B(n2647), .Y(n1196) );
  OAI21X1TS U690 ( .A0(n1250), .A1(n2647), .B0(n1196), .Y(n971) );
  NAND2X1TS U691 ( .A(n1487), .B(n1513), .Y(\DP_OP_159_297_3515/n1014 ) );
  XNOR2X4TS U692 ( .A(n1199), .B(n1200), .Y(n1198) );
  INVX12TS U693 ( .A(\add_x_22_4/n30 ), .Y(n1200) );
  NOR2BX4TS U694 ( .AN(\add_x_22_4/n34 ), .B(n1201), .Y(n1199) );
  INVX12TS U695 ( .A(n2031), .Y(n1201) );
  NAND2BX1TS U696 ( .AN(n1198), .B(n1713), .Y(n1197) );
  OAI2BB1X1TS U697 ( .A0N(n2565), .A1N(n2653), .B0(n1197), .Y(n948) );
  XNOR2X4TS U698 ( .A(n1204), .B(n1205), .Y(n1203) );
  INVX12TS U699 ( .A(\add_x_22_2/n12 ), .Y(n1205) );
  NOR2BX4TS U700 ( .AN(\add_x_22_2/n16 ), .B(n1206), .Y(n1204) );
  INVX12TS U701 ( .A(n2582), .Y(n1206) );
  NAND2X1TS U702 ( .A(n1724), .B(\addr_calc/fft_write_calc/counter/N61 ), .Y(
        n1207) );
  OAI2BB1X2TS U703 ( .A0N(\addr_calc/fft_write_calc/count[18] ), .A1N(n2664), 
        .B0(n1207), .Y(n1048) );
  NOR2X4TS U704 ( .A(n1795), .B(\DP_OP_158_296_6262/n1889 ), .Y(
        \DP_OP_158_296_6262/n1888 ) );
  XNOR2X4TS U705 ( .A(\DP_OP_158_296_6262/n1888 ), .B(n1516), .Y(n1652) );
  XNOR2X1TS U706 ( .A(n2372), .B(\addr_calc/fft_write_calc/count[0] ), .Y(
        \DP_OP_158_296_6262/n822 ) );
  XOR2X1TS U707 ( .A(n2596), .B(n2032), .Y(n1208) );
  XOR2X1TS U708 ( .A(\DP_OP_158_296_6262/n855 ), .B(
        \addr_calc/fft_write_calc/count[4] ), .Y(n1211) );
  XOR2X1TS U709 ( .A(n2599), .B(n2568), .Y(n1210) );
  XOR2X1TS U710 ( .A(n2593), .B(n2030), .Y(n1209) );
  XOR2X1TS U711 ( .A(n2595), .B(n1479), .Y(n1212) );
  XOR2X4TS U712 ( .A(n1777), .B(n1852), .Y(\DP_OP_158_296_6262/n486 ) );
  XNOR2X4TS U713 ( .A(n1718), .B(n2011), .Y(\DP_OP_158_296_6262/n566 ) );
  XOR2X4TS U714 ( .A(n1655), .B(n1915), .Y(n1213) );
  XNOR2X2TS U715 ( .A(n2602), .B(n1913), .Y(\DP_OP_158_296_6262/n515 ) );
  XNOR2X2TS U716 ( .A(n1652), .B(n2014), .Y(\DP_OP_158_296_6262/n595 ) );
  XNOR2X1TS U717 ( .A(\DP_OP_158_296_6262/n838 ), .B(n1918), .Y(
        \DP_OP_158_296_6262/n608 ) );
  XNOR2X1TS U718 ( .A(n1660), .B(n1667), .Y(\DP_OP_158_296_6262/n733 ) );
  XNOR2X1TS U719 ( .A(n1976), .B(n1658), .Y(\DP_OP_158_296_6262/n689 ) );
  XNOR2X2TS U720 ( .A(n1657), .B(n2021), .Y(\DP_OP_158_296_6262/n702 ) );
  XNOR2X2TS U721 ( .A(n1729), .B(\addr_calc/fft_write_calc/count[17] ), .Y(
        \DP_OP_158_296_6262/n664 ) );
  XOR2X4TS U722 ( .A(\DP_OP_158_296_6262/n841 ), .B(n2019), .Y(
        \DP_OP_158_296_6262/n649 ) );
  XNOR2X2TS U723 ( .A(n1654), .B(n1922), .Y(\DP_OP_158_296_6262/n632 ) );
  XOR2X2TS U724 ( .A(\DP_OP_158_296_6262/n829 ), .B(n1849), .Y(n1216) );
  NOR2X2TS U725 ( .A(\DP_OP_158_296_6262/n501 ), .B(\DP_OP_158_296_6262/n486 ), 
        .Y(\DP_OP_158_296_6262/n484 ) );
  NOR2BX4TS U726 ( .AN(n1213), .B(\DP_OP_158_296_6262/n566 ), .Y(
        \DP_OP_158_296_6262/n549 ) );
  NOR2X2TS U727 ( .A(\DP_OP_158_296_6262/n595 ), .B(\DP_OP_158_296_6262/n580 ), 
        .Y(\DP_OP_158_296_6262/n578 ) );
  NOR2X2TS U728 ( .A(\DP_OP_158_296_6262/n621 ), .B(\DP_OP_158_296_6262/n608 ), 
        .Y(\DP_OP_158_296_6262/n606 ) );
  NOR2X2TS U729 ( .A(\DP_OP_158_296_6262/n769 ), .B(\DP_OP_158_296_6262/n776 ), 
        .Y(\DP_OP_158_296_6262/n767 ) );
  NOR2X1TS U730 ( .A(\DP_OP_158_296_6262/n753 ), .B(\DP_OP_158_296_6262/n762 ), 
        .Y(\DP_OP_158_296_6262/n751 ) );
  NOR2X2TS U731 ( .A(\DP_OP_158_296_6262/n744 ), .B(\DP_OP_158_296_6262/n733 ), 
        .Y(\DP_OP_158_296_6262/n731 ) );
  NOR2X2TS U732 ( .A(\DP_OP_158_296_6262/n724 ), .B(\DP_OP_158_296_6262/n713 ), 
        .Y(\DP_OP_158_296_6262/n711 ) );
  NOR2X2TS U733 ( .A(\DP_OP_158_296_6262/n664 ), .B(\DP_OP_158_296_6262/n677 ), 
        .Y(\DP_OP_158_296_6262/n662 ) );
  NOR2X2TS U734 ( .A(\DP_OP_158_296_6262/n632 ), .B(\DP_OP_158_296_6262/n649 ), 
        .Y(\DP_OP_158_296_6262/n630 ) );
  NAND2X2TS U735 ( .A(\DP_OP_158_296_6262/n484 ), .B(n1216), .Y(
        \DP_OP_158_296_6262/n465 ) );
  NAND2X4TS U736 ( .A(\DP_OP_158_296_6262/n513 ), .B(\DP_OP_158_296_6262/n549 ), .Y(\DP_OP_158_296_6262/n511 ) );
  NAND2X1TS U737 ( .A(\DP_OP_158_296_6262/n731 ), .B(\DP_OP_158_296_6262/n751 ), .Y(\DP_OP_158_296_6262/n729 ) );
  NAND2X2TS U738 ( .A(\DP_OP_158_296_6262/n687 ), .B(\DP_OP_158_296_6262/n711 ), .Y(\DP_OP_158_296_6262/n685 ) );
  NAND2X2TS U739 ( .A(\DP_OP_158_296_6262/n630 ), .B(\DP_OP_158_296_6262/n662 ), .Y(\DP_OP_158_296_6262/n628 ) );
  NOR2X2TS U740 ( .A(\DP_OP_158_296_6262/n465 ), .B(\DP_OP_158_296_6262/n452 ), 
        .Y(\DP_OP_158_296_6262/n450 ) );
  NOR2X4TS U741 ( .A(\DP_OP_158_296_6262/n576 ), .B(\DP_OP_158_296_6262/n511 ), 
        .Y(\DP_OP_158_296_6262/n509 ) );
  AND2X8TS U742 ( .A(\DP_OP_158_296_6262/n509 ), .B(\DP_OP_158_296_6262/n450 ), 
        .Y(n1214) );
  AND2X8TS U743 ( .A(\DP_OP_158_296_6262/n626 ), .B(\DP_OP_158_296_6262/n727 ), 
        .Y(n1215) );
  NAND2X8TS U744 ( .A(n1215), .B(n1214), .Y(
        \addr_calc/fft_write_calc/counter/N38 ) );
  AOI21X4TS U745 ( .A0(\addr_calc/fft_write_calc/counter/N38 ), .A1(
        data_from_fft), .B0(n2586), .Y(n2797) );
  NAND2BX4TS U746 ( .AN(n1218), .B(n1724), .Y(n1217) );
  XNOR2X4TS U747 ( .A(\add_x_22_1/n34 ), .B(n1219), .Y(n1218) );
  INVX12TS U748 ( .A(n2013), .Y(n1219) );
  OAI2BB1X2TS U749 ( .A0N(\addr_calc/fft_write_calc/count[22] ), .A1N(n2667), 
        .B0(n1217), .Y(n1044) );
  XNOR2X4TS U750 ( .A(\add_x_22_1/n41 ), .B(n1222), .Y(n1221) );
  INVX12TS U751 ( .A(n2016), .Y(n1222) );
  NAND2BX1TS U752 ( .AN(n1221), .B(n1722), .Y(n1220) );
  OAI2BB1X2TS U753 ( .A0N(\addr_calc/fft_write_calc/count[20] ), .A1N(n2666), 
        .B0(n1220), .Y(n1046) );
  INVX12TS U754 ( .A(n1616), .Y(n1223) );
  NAND2BX1TS U755 ( .AN(n1758), .B(\addr_calc/fir_write_calc/counter/N53 ), 
        .Y(n1226) );
  OAI2BB1X1TS U756 ( .A0N(n1874), .A1N(n1263), .B0(n1226), .Y(n1120) );
  NAND2BX1TS U757 ( .AN(n1758), .B(\addr_calc/fir_write_calc/counter/N50 ), 
        .Y(n1225) );
  OAI2BB1X1TS U758 ( .A0N(n1869), .A1N(n1269), .B0(n1225), .Y(n1123) );
  NAND2BX1TS U759 ( .AN(n1758), .B(\addr_calc/fir_write_calc/counter/N44 ), 
        .Y(n1224) );
  OAI2BB1X1TS U760 ( .A0N(n1868), .A1N(n1261), .B0(n1224), .Y(n1129) );
  NAND2BX1TS U761 ( .AN(n1758), .B(n1223), .Y(n1615) );
  OAI2BB1X4TS U762 ( .A0N(\add_x_19_2/n59 ), .A1N(n1231), .B0(n1232), .Y(n1230) );
  OAI2BB1X4TS U763 ( .A0N(\add_x_19_2/n58 ), .A1N(\add_x_19_2/n59 ), .B0(n1233), .Y(n1232) );
  INVX12TS U764 ( .A(n1231), .Y(n1233) );
  NOR2BX4TS U765 ( .AN(\add_x_19_2/n59 ), .B(n1231), .Y(n1229) );
  NAND2BX4TS U766 ( .AN(\add_x_19_2/n58 ), .B(n1231), .Y(n1227) );
  NOR2BX4TS U767 ( .AN(\add_x_19_2/n56 ), .B(\add_x_19_2/n55 ), .Y(n1231) );
  NOR2X4TS U768 ( .A(n1493), .B(n1497), .Y(\DP_OP_158_296_6262/n1999 ) );
  NOR2X2TS U769 ( .A(n1495), .B(n1489), .Y(\DP_OP_158_296_6262/n1988 ) );
  NAND2X4TS U770 ( .A(\DP_OP_158_296_6262/n1999 ), .B(
        \DP_OP_158_296_6262/n1988 ), .Y(\DP_OP_158_296_6262/n1987 ) );
  NOR2BX4TS U771 ( .AN(n1641), .B(n1527), .Y(n1234) );
  NAND2X6TS U772 ( .A(n1797), .B(n1234), .Y(\DP_OP_158_296_6262/n2011 ) );
  NAND2X2TS U773 ( .A(\DP_OP_158_296_6262/n1945 ), .B(
        \DP_OP_158_296_6262/n1933 ), .Y(\DP_OP_158_296_6262/n1932 ) );
  NOR2X4TS U774 ( .A(\DP_OP_158_296_6262/n1958 ), .B(
        \DP_OP_158_296_6262/n1932 ), .Y(\DP_OP_158_296_6262/n1931 ) );
  NOR2X4TS U775 ( .A(n1795), .B(n2361), .Y(\DP_OP_158_296_6262/n1923 ) );
  XNOR2X4TS U776 ( .A(\DP_OP_158_296_6262/n1923 ), .B(n2369), .Y(n1729) );
  XNOR2X1TS U777 ( .A(n2372), .B(n1986), .Y(\DP_OP_158_296_6262/n1716 ) );
  XOR2X1TS U778 ( .A(n2596), .B(\addr_calc/fir_write_calc/count[2] ), .Y(n1235) );
  XOR2X1TS U779 ( .A(\DP_OP_158_296_6262/n855 ), .B(n1865), .Y(n1238) );
  XOR2X1TS U780 ( .A(n2599), .B(n1866), .Y(n1237) );
  XOR2X1TS U781 ( .A(n2593), .B(n1992), .Y(n1236) );
  XOR2X1TS U782 ( .A(n2595), .B(\addr_calc/fir_write_calc/count[5] ), .Y(n1239) );
  XNOR2X1TS U783 ( .A(n1872), .B(n1469), .Y(\DP_OP_158_296_6262/n1647 ) );
  XNOR2X1TS U784 ( .A(n1874), .B(n1656), .Y(\DP_OP_158_296_6262/n1638 ) );
  XNOR2X1TS U785 ( .A(n1880), .B(n1659), .Y(\DP_OP_158_296_6262/n1607 ) );
  XNOR2X2TS U786 ( .A(n1756), .B(n1999), .Y(\DP_OP_158_296_6262/n1618 ) );
  XNOR2X2TS U787 ( .A(n1729), .B(n1886), .Y(\DP_OP_158_296_6262/n1558 ) );
  XNOR2X4TS U788 ( .A(\DP_OP_158_296_6262/n841 ), .B(
        \addr_calc/fir_write_calc/count[18] ), .Y(\DP_OP_158_296_6262/n1543 )
         );
  XNOR2X2TS U789 ( .A(n1654), .B(\addr_calc/fir_write_calc/count[19] ), .Y(
        \DP_OP_158_296_6262/n1526 ) );
  XNOR2X4TS U790 ( .A(n1463), .B(\addr_calc/fir_write_calc/count[29] ), .Y(
        \DP_OP_158_296_6262/n1380 ) );
  XOR2X4TS U791 ( .A(n1718), .B(\add_x_22_3/n22 ), .Y(
        \DP_OP_158_296_6262/n1460 ) );
  XNOR2X2TS U792 ( .A(n1655), .B(n1894), .Y(\DP_OP_158_296_6262/n1445 ) );
  XNOR2X2TS U793 ( .A(n2602), .B(\addr_calc/fir_write_calc/count[27] ), .Y(
        \DP_OP_158_296_6262/n1409 ) );
  XNOR2X4TS U794 ( .A(\DP_OP_158_296_6262/n833 ), .B(n2581), .Y(
        \DP_OP_158_296_6262/n1428 ) );
  XOR2X2TS U795 ( .A(\DP_OP_158_296_6262/n838 ), .B(n1891), .Y(
        \DP_OP_158_296_6262/n1502 ) );
  XNOR2X2TS U796 ( .A(n1776), .B(n2009), .Y(\DP_OP_158_296_6262/n1515 ) );
  XNOR2X4TS U797 ( .A(n1730), .B(n2563), .Y(\DP_OP_158_296_6262/n1474 ) );
  XNOR2X2TS U798 ( .A(n1652), .B(\addr_calc/fir_write_calc/count[22] ), .Y(
        \DP_OP_158_296_6262/n1489 ) );
  NOR2X2TS U799 ( .A(\DP_OP_158_296_6262/n1663 ), .B(
        \DP_OP_158_296_6262/n1670 ), .Y(\DP_OP_158_296_6262/n1661 ) );
  NOR2X2TS U800 ( .A(\DP_OP_158_296_6262/n1647 ), .B(
        \DP_OP_158_296_6262/n1656 ), .Y(\DP_OP_158_296_6262/n1645 ) );
  NOR2X2TS U801 ( .A(\DP_OP_158_296_6262/n1638 ), .B(
        \DP_OP_158_296_6262/n1627 ), .Y(\DP_OP_158_296_6262/n1625 ) );
  NOR2X2TS U802 ( .A(\DP_OP_158_296_6262/n1596 ), .B(
        \DP_OP_158_296_6262/n1583 ), .Y(\DP_OP_158_296_6262/n1581 ) );
  NOR2X2TS U803 ( .A(\DP_OP_158_296_6262/n1618 ), .B(
        \DP_OP_158_296_6262/n1607 ), .Y(\DP_OP_158_296_6262/n1605 ) );
  NOR2X4TS U804 ( .A(\DP_OP_158_296_6262/n1558 ), .B(
        \DP_OP_158_296_6262/n1571 ), .Y(\DP_OP_158_296_6262/n1556 ) );
  NOR2X4TS U805 ( .A(\DP_OP_158_296_6262/n1526 ), .B(
        \DP_OP_158_296_6262/n1543 ), .Y(\DP_OP_158_296_6262/n1524 ) );
  XOR2X2TS U806 ( .A(\DP_OP_158_296_6262/n829 ), .B(
        \addr_calc/fir_write_calc/count[30] ), .Y(n1240) );
  NOR2X2TS U807 ( .A(\DP_OP_158_296_6262/n1380 ), .B(
        \DP_OP_158_296_6262/n1395 ), .Y(\DP_OP_158_296_6262/n1378 ) );
  NOR2X4TS U808 ( .A(\DP_OP_158_296_6262/n1445 ), .B(
        \DP_OP_158_296_6262/n1460 ), .Y(\DP_OP_158_296_6262/n1443 ) );
  NOR2X4TS U809 ( .A(\DP_OP_158_296_6262/n1428 ), .B(
        \DP_OP_158_296_6262/n1409 ), .Y(\DP_OP_158_296_6262/n1407 ) );
  NOR2X2TS U810 ( .A(\DP_OP_158_296_6262/n1515 ), .B(
        \DP_OP_158_296_6262/n1502 ), .Y(\DP_OP_158_296_6262/n1500 ) );
  NOR2X2TS U811 ( .A(\DP_OP_158_296_6262/n1489 ), .B(
        \DP_OP_158_296_6262/n1474 ), .Y(\DP_OP_158_296_6262/n1472 ) );
  NAND2X2TS U812 ( .A(\DP_OP_158_296_6262/n1661 ), .B(
        \DP_OP_158_296_6262/n1688 ), .Y(\DP_OP_158_296_6262/n1659 ) );
  NAND2X2TS U813 ( .A(\DP_OP_158_296_6262/n1625 ), .B(
        \DP_OP_158_296_6262/n1645 ), .Y(\DP_OP_158_296_6262/n1623 ) );
  NAND2X2TS U814 ( .A(\DP_OP_158_296_6262/n1605 ), .B(
        \DP_OP_158_296_6262/n1581 ), .Y(\DP_OP_158_296_6262/n1579 ) );
  NAND2X4TS U815 ( .A(\DP_OP_158_296_6262/n1524 ), .B(
        \DP_OP_158_296_6262/n1556 ), .Y(\DP_OP_158_296_6262/n1522 ) );
  NAND2X2TS U816 ( .A(\DP_OP_158_296_6262/n1378 ), .B(n1240), .Y(
        \DP_OP_158_296_6262/n1359 ) );
  NAND2X4TS U817 ( .A(\DP_OP_158_296_6262/n1407 ), .B(
        \DP_OP_158_296_6262/n1443 ), .Y(\DP_OP_158_296_6262/n1405 ) );
  NAND2X2TS U818 ( .A(\DP_OP_158_296_6262/n1472 ), .B(
        \DP_OP_158_296_6262/n1500 ), .Y(\DP_OP_158_296_6262/n1470 ) );
  NOR2X4TS U819 ( .A(\DP_OP_158_296_6262/n1623 ), .B(
        \DP_OP_158_296_6262/n1659 ), .Y(\DP_OP_158_296_6262/n1621 ) );
  NOR2X4TS U820 ( .A(\DP_OP_158_296_6262/n1522 ), .B(
        \DP_OP_158_296_6262/n1579 ), .Y(\DP_OP_158_296_6262/n1520 ) );
  NOR2X2TS U821 ( .A(\DP_OP_158_296_6262/n1359 ), .B(
        \DP_OP_158_296_6262/n1346 ), .Y(\DP_OP_158_296_6262/n1344 ) );
  NOR2X4TS U822 ( .A(\DP_OP_158_296_6262/n1470 ), .B(
        \DP_OP_158_296_6262/n1405 ), .Y(\DP_OP_158_296_6262/n1403 ) );
  NAND2X4TS U823 ( .A(\DP_OP_158_296_6262/n1520 ), .B(
        \DP_OP_158_296_6262/n1621 ), .Y(\DP_OP_158_296_6262/n1518 ) );
  NAND2X2TS U824 ( .A(\DP_OP_158_296_6262/n1403 ), .B(
        \DP_OP_158_296_6262/n1344 ), .Y(\DP_OP_158_296_6262/n1342 ) );
  OR2X8TS U825 ( .A(\DP_OP_158_296_6262/n1342 ), .B(\DP_OP_158_296_6262/n1518 ), .Y(\addr_calc/fir_write_calc/counter/N38 ) );
  OR3X1TS U826 ( .A(\data_cntl/N95 ), .B(n2804), .C(n2061), .Y(n1241) );
  CLKINVX1TS U827 ( .A(n1868), .Y(\add_x_22_3/n121 ) );
  XNOR2X1TS U828 ( .A(\add_x_22_3/n121 ), .B(
        \addr_calc/fir_write_calc/count[0] ), .Y(
        \addr_calc/fir_write_calc/counter/N44 ) );
  XNOR2X4TS U829 ( .A(\add_x_22_1/n102 ), .B(n1244), .Y(n1243) );
  INVX12TS U830 ( .A(n2029), .Y(n1244) );
  NAND2BX1TS U831 ( .AN(n1243), .B(n1145), .Y(n1242) );
  OAI2BB1X1TS U832 ( .A0N(\addr_calc/fft_write_calc/count[6] ), .A1N(n2663), 
        .B0(n1242), .Y(n1060) );
  NAND2X2TS U833 ( .A(\DP_OP_159_297_3515/n1064 ), .B(
        \DP_OP_159_297_3515/n1040 ), .Y(\DP_OP_159_297_3515/n1039 ) );
  NOR2X1TS U834 ( .A(\DP_OP_159_297_3515/n998 ), .B(\DP_OP_159_297_3515/n986 ), 
        .Y(\DP_OP_159_297_3515/n985 ) );
  AND2X4TS U835 ( .A(\DP_OP_159_297_3515/n985 ), .B(\DP_OP_159_297_3515/n1011 ), .Y(n1245) );
  NAND2BX4TS U836 ( .AN(\DP_OP_159_297_3515/n1039 ), .B(n1245), .Y(n1782) );
  CLKINVX1TS U837 ( .A(\DP_OP_159_297_3515/n971 ), .Y(
        \DP_OP_159_297_3515/n970 ) );
  NAND2X2TS U838 ( .A(n1790), .B(\DP_OP_159_297_3515/n970 ), .Y(
        \DP_OP_159_297_3515/n969 ) );
  XNOR2X4TS U839 ( .A(\DP_OP_159_297_3515/n969 ), .B(\DP_OP_159_297_3515/n964 ), .Y(n1662) );
  XNOR2X1TS U840 ( .A(\addr_calc/iir_read_calc/count[0] ), .B(
        \DP_OP_159_297_3515/n815 ), .Y(\DP_OP_159_297_3515/n353 ) );
  XOR2X1TS U841 ( .A(n2612), .B(\addr_calc/iir_read_calc/count[2] ), .Y(n1246)
         );
  XOR2X1TS U842 ( .A(n2624), .B(n1903), .Y(n1248) );
  NOR2X2TS U843 ( .A(\DP_OP_159_297_3515/n343 ), .B(\DP_OP_159_297_3515/n341 ), 
        .Y(\DP_OP_159_297_3515/n339 ) );
  XOR2X1TS U844 ( .A(n2623), .B(n2553), .Y(n1249) );
  XOR2X1TS U845 ( .A(n2610), .B(n2018), .Y(n1247) );
  NAND2X2TS U846 ( .A(\DP_OP_159_297_3515/n339 ), .B(n1248), .Y(
        \DP_OP_159_297_3515/n333 ) );
  XNOR2X2TS U847 ( .A(n2622), .B(n2583), .Y(\DP_OP_159_297_3515/n305 ) );
  XNOR2X1TS U848 ( .A(n2608), .B(\addr_calc/iir_read_calc/count[9] ), .Y(
        \DP_OP_159_297_3515/n298 ) );
  XNOR2X2TS U849 ( .A(n2620), .B(\addr_calc/iir_read_calc/count[11] ), .Y(
        \DP_OP_159_297_3515/n280 ) );
  XOR2X4TS U850 ( .A(n2618), .B(\add_x_22_4/n71 ), .Y(
        \DP_OP_159_297_3515/n260 ) );
  XNOR2X4TS U851 ( .A(n2617), .B(n1784), .Y(\DP_OP_159_297_3515/n249 ) );
  XNOR2X4TS U852 ( .A(n2615), .B(n1916), .Y(\DP_OP_159_297_3515/n225 ) );
  XNOR2X4TS U853 ( .A(n2616), .B(n2566), .Y(\DP_OP_159_297_3515/n238 ) );
  XNOR2X4TS U854 ( .A(\DP_OP_159_297_3515/n1128 ), .B(n2024), .Y(
        \DP_OP_159_297_3515/n200 ) );
  XNOR2X2TS U855 ( .A(n2607), .B(\addr_calc/iir_read_calc/count[17] ), .Y(
        \DP_OP_159_297_3515/n213 ) );
  XNOR2X4TS U856 ( .A(n1662), .B(n2556), .Y(\DP_OP_159_297_3515/n185 ) );
  XOR2X4TS U857 ( .A(n1697), .B(n2027), .Y(\DP_OP_159_297_3515/n168 ) );
  NOR2X2TS U858 ( .A(\DP_OP_159_297_3515/n317 ), .B(\DP_OP_159_297_3515/n333 ), 
        .Y(\DP_OP_159_297_3515/n315 ) );
  NOR2X2TS U859 ( .A(\DP_OP_159_297_3515/n305 ), .B(\DP_OP_159_297_3515/n312 ), 
        .Y(\DP_OP_159_297_3515/n303 ) );
  NOR2X4TS U860 ( .A(\DP_OP_159_297_3515/n289 ), .B(\DP_OP_159_297_3515/n298 ), 
        .Y(\DP_OP_159_297_3515/n287 ) );
  NOR2X4TS U861 ( .A(\DP_OP_159_297_3515/n280 ), .B(\DP_OP_159_297_3515/n269 ), 
        .Y(\DP_OP_159_297_3515/n267 ) );
  NOR2X4TS U862 ( .A(\DP_OP_159_297_3515/n249 ), .B(\DP_OP_159_297_3515/n260 ), 
        .Y(\DP_OP_159_297_3515/n247 ) );
  NOR2X4TS U863 ( .A(\DP_OP_159_297_3515/n238 ), .B(\DP_OP_159_297_3515/n225 ), 
        .Y(\DP_OP_159_297_3515/n223 ) );
  NOR2X4TS U864 ( .A(\DP_OP_159_297_3515/n213 ), .B(\DP_OP_159_297_3515/n200 ), 
        .Y(\DP_OP_159_297_3515/n198 ) );
  NOR2X8TS U865 ( .A(\DP_OP_159_297_3515/n168 ), .B(\DP_OP_159_297_3515/n185 ), 
        .Y(\DP_OP_159_297_3515/n166 ) );
  NAND2X2TS U866 ( .A(\DP_OP_159_297_3515/n303 ), .B(\DP_OP_159_297_3515/n315 ), .Y(\DP_OP_159_297_3515/n301 ) );
  NAND2X4TS U867 ( .A(\DP_OP_159_297_3515/n267 ), .B(\DP_OP_159_297_3515/n287 ), .Y(\DP_OP_159_297_3515/n265 ) );
  NAND2X2TS U868 ( .A(\DP_OP_159_297_3515/n223 ), .B(\DP_OP_159_297_3515/n247 ), .Y(\DP_OP_159_297_3515/n221 ) );
  NAND2X4TS U869 ( .A(\DP_OP_159_297_3515/n166 ), .B(\DP_OP_159_297_3515/n198 ), .Y(\DP_OP_159_297_3515/n164 ) );
  NOR2X4TS U870 ( .A(\DP_OP_159_297_3515/n265 ), .B(\DP_OP_159_297_3515/n301 ), 
        .Y(\DP_OP_159_297_3515/n263 ) );
  NOR2X4TS U871 ( .A(\DP_OP_159_297_3515/n164 ), .B(\DP_OP_159_297_3515/n221 ), 
        .Y(\DP_OP_159_297_3515/n162 ) );
  NAND2X4TS U872 ( .A(\DP_OP_159_297_3515/n162 ), .B(\DP_OP_159_297_3515/n263 ), .Y(\DP_OP_159_297_3515/n160 ) );
  OR2X8TS U873 ( .A(\DP_OP_159_297_3515/n1 ), .B(\DP_OP_159_297_3515/n160 ), 
        .Y(\addr_calc/iir_read_calc/counter/N38 ) );
  OAI21XLTS U874 ( .A0(n2786), .A1(n2785), .B0(iir_enable), .Y(n1250) );
  XNOR2X4TS U875 ( .A(n1254), .B(\add_x_22_4/n71 ), .Y(n1253) );
  NAND2BX4TS U876 ( .AN(n1255), .B(\add_x_22_4/n75 ), .Y(n1254) );
  INVX12TS U877 ( .A(n1785), .Y(n1255) );
  INVX12TS U878 ( .A(\add_x_22_4/n71 ), .Y(n1251) );
  NAND2BX1TS U879 ( .AN(n1253), .B(n1713), .Y(n1252) );
  OAI2BB1X2TS U880 ( .A0N(n1251), .A1N(n2649), .B0(n1252), .Y(n958) );
  NOR2X4TS U881 ( .A(\DP_OP_158_296_6262/n1176 ), .B(
        \DP_OP_158_296_6262/n1212 ), .Y(\DP_OP_158_296_6262/n1174 ) );
  INVX3TS U882 ( .A(n2805), .Y(n1256) );
  INVX2TS U883 ( .A(n2805), .Y(n1257) );
  INVX2TS U884 ( .A(n2805), .Y(n1258) );
  INVX3TS U885 ( .A(n1256), .Y(n1259) );
  CLKINVX3TS U886 ( .A(n1256), .Y(n1260) );
  CLKINVX3TS U887 ( .A(n1256), .Y(n1261) );
  CLKINVX3TS U888 ( .A(n1256), .Y(n1262) );
  CLKINVX3TS U889 ( .A(n1257), .Y(n1263) );
  CLKINVX3TS U890 ( .A(n1257), .Y(n1264) );
  CLKINVX3TS U891 ( .A(n1257), .Y(n1265) );
  CLKINVX3TS U892 ( .A(n1257), .Y(n1266) );
  CLKINVX3TS U893 ( .A(n1258), .Y(n1267) );
  CLKINVX3TS U894 ( .A(n1258), .Y(n1268) );
  CLKINVX3TS U895 ( .A(n1258), .Y(n1269) );
  CLKINVX3TS U896 ( .A(n1258), .Y(n1270) );
  OAI2BB1X2TS U897 ( .A0N(n1865), .A1N(n1266), .B0(n1615), .Y(n1126) );
  XOR2X4TS U898 ( .A(n2625), .B(n1684), .Y(n1623) );
  XNOR2X2TS U899 ( .A(n2614), .B(\addr_calc/iir_write_calc/count[31] ), .Y(
        \DP_OP_159_297_3515/n430 ) );
  CLKINVX3TS U900 ( .A(\DP_OP_159_297_3515/n1024 ), .Y(n1733) );
  XNOR2X2TS U901 ( .A(n2613), .B(n1850), .Y(n1563) );
  XOR2X2TS U902 ( .A(n1693), .B(n2364), .Y(n2598) );
  NOR2X1TS U903 ( .A(\add_x_19_5/n123 ), .B(\add_x_19_5/n120 ), .Y(
        \add_x_19_5/n118 ) );
  NOR2X1TS U904 ( .A(n1944), .B(n2500), .Y(\add_x_19_0/n55 ) );
  NOR2X1TS U905 ( .A(n1688), .B(n2498), .Y(\add_x_19_5/n55 ) );
  OR4X6TS U906 ( .A(n783), .B(n2793), .C(\data_cntl/N63 ), .D(n2588), .Y(n1701) );
  NOR2X1TS U907 ( .A(n1879), .B(n2450), .Y(\add_x_19_2/n86 ) );
  NOR2X1TS U908 ( .A(n1556), .B(n1557), .Y(n1555) );
  NOR2X1TS U909 ( .A(n1845), .B(n2380), .Y(n1557) );
  AND2X2TS U910 ( .A(\addr_calc/fft_write_calc/count[31] ), .B(n2380), .Y(
        n1556) );
  NOR2BX1TS U911 ( .AN(\add_x_19_1/n37 ), .B(n1555), .Y(n1552) );
  INVX2TS U912 ( .A(n1555), .Y(n1554) );
  INVX2TS U913 ( .A(\add_x_19_1/n42 ), .Y(n1546) );
  NOR2BX1TS U914 ( .AN(\add_x_22_5/n68 ), .B(\add_x_22_5/n67 ), .Y(n1575) );
  NOR2BX1TS U915 ( .AN(\add_x_22_4/n16 ), .B(\add_x_22_4/n15 ), .Y(n1578) );
  NOR2BX1TS U916 ( .AN(n1972), .B(\add_x_22_0/n85 ), .Y(n1622) );
  INVX2TS U917 ( .A(\add_x_22_0/n101 ), .Y(n1610) );
  INVX2TS U918 ( .A(\add_x_22_4/n15 ), .Y(n1572) );
  AOI21X2TS U919 ( .A0(\add_x_19_0/n43 ), .A1(n2628), .B0(n1541), .Y(
        \add_x_19_0/n38 ) );
  INVX2TS U920 ( .A(\add_x_19_0/n42 ), .Y(n1541) );
  NOR2X1TS U921 ( .A(n1835), .B(n2500), .Y(\add_x_19_3/n55 ) );
  INVX2TS U922 ( .A(\add_x_19_3/n42 ), .Y(n1535) );
  NOR2BX1TS U923 ( .AN(\add_x_19_5/n59 ), .B(n1607), .Y(n1605) );
  NOR2BX1TS U924 ( .AN(\add_x_19_5/n56 ), .B(\add_x_19_5/n55 ), .Y(n1607) );
  NOR2BX1TS U925 ( .AN(n2554), .B(\add_x_22_0/n58 ), .Y(n1635) );
  NAND2BX1TS U926 ( .AN(\add_x_22_0/n40 ), .B(\add_x_22_0/n41 ), .Y(n1629) );
  INVX4TS U927 ( .A(n1701), .Y(n1752) );
  INVX2TS U928 ( .A(\addr_calc/iir_read_calc/count[26] ), .Y(\add_x_22_4/n15 )
         );
  XNOR2X1TS U929 ( .A(\DP_OP_158_296_6262/n2015 ), .B(n2363), .Y(n2599) );
  NOR2X1TS U930 ( .A(\add_x_19_2/n123 ), .B(\add_x_19_2/n120 ), .Y(
        \add_x_19_2/n118 ) );
  XNOR2X1TS U931 ( .A(\DP_OP_158_296_6262/n838 ), .B(
        \addr_calc/fir_read_calc/count[21] ), .Y(\DP_OP_158_296_6262/n161 ) );
  NOR2BX1TS U932 ( .AN(n1626), .B(n2796), .Y(n1625) );
  NOR2X1TS U933 ( .A(n2587), .B(\data_cntl/N9 ), .Y(n1626) );
  OAI21X1TS U934 ( .A0(\add_x_19_3/n120 ), .A1(\add_x_19_3/n124 ), .B0(
        \add_x_19_3/n121 ), .Y(n1595) );
  NOR2X1TS U935 ( .A(\add_x_19_0/n162 ), .B(\add_x_19_0/n165 ), .Y(n1558) );
  INVX2TS U936 ( .A(n1491), .Y(\DP_OP_158_296_6262/n1897 ) );
  NOR2X1TS U937 ( .A(n1926), .B(n2492), .Y(\add_x_19_4/n63 ) );
  NOR2X1TS U938 ( .A(n1950), .B(n2469), .Y(\add_x_19_0/n78 ) );
  OAI21X1TS U939 ( .A0(\add_x_19_0/n90 ), .A1(\add_x_19_0/n86 ), .B0(
        \add_x_19_0/n87 ), .Y(\add_x_19_0/n85 ) );
  NOR2X1TS U940 ( .A(\DP_OP_158_296_6262/n306 ), .B(\DP_OP_158_296_6262/n315 ), 
        .Y(\DP_OP_158_296_6262/n304 ) );
  NOR2X1TS U941 ( .A(n1689), .B(n2475), .Y(\add_x_19_0/n120 ) );
  NOR2X1TS U942 ( .A(n1965), .B(n2470), .Y(\add_x_19_5/n78 ) );
  NOR4XLTS U943 ( .A(\addr_calc/iir_write_calc/count[30] ), .B(n2036), .C(
        \addr_calc/iir_write_calc/count[29] ), .D(n1974), .Y(n918) );
  NOR2X1TS U944 ( .A(\add_x_19_4/n66 ), .B(\add_x_19_4/n63 ), .Y(
        \add_x_19_4/n61 ) );
  NOR2X1TS U945 ( .A(n1913), .B(n2498), .Y(\add_x_19_1/n55 ) );
  CLKINVX6TS U946 ( .A(n2813), .Y(n1765) );
  NOR2X1TS U947 ( .A(n1667), .B(n2404), .Y(\add_x_19_1/n139 ) );
  NOR2X1TS U948 ( .A(\add_x_19_5/n135 ), .B(\add_x_19_5/n116 ), .Y(
        \add_x_19_5/n114 ) );
  NOR2X1TS U949 ( .A(n2384), .B(n1871), .Y(\add_x_19_2/n48 ) );
  OAI21XLTS U950 ( .A0(\add_x_19_0/n181 ), .A1(\add_x_19_0/n185 ), .B0(
        \add_x_19_0/n182 ), .Y(n1588) );
  OAI21X1TS U951 ( .A0(\add_x_19_2/n181 ), .A1(\add_x_19_2/n185 ), .B0(
        \add_x_19_2/n182 ), .Y(n1548) );
  OAI21X1TS U952 ( .A0(\add_x_19_1/n191 ), .A1(\add_x_19_1/n188 ), .B0(
        \add_x_19_1/n189 ), .Y(\add_x_19_1/n187 ) );
  INVX2TS U953 ( .A(n2065), .Y(n2066) );
  CLKBUFX2TS U954 ( .A(n2074), .Y(n2584) );
  INVX2TS U955 ( .A(n1494), .Y(n1495) );
  NOR2X1TS U956 ( .A(n2021), .B(n2425), .Y(\add_x_19_1/n123 ) );
  NOR2X1TS U957 ( .A(n1958), .B(n2487), .Y(\add_x_19_5/n97 ) );
  INVXLTS U958 ( .A(\addr_calc/iir_read_calc/count[14] ), .Y(\add_x_22_4/n67 )
         );
  INVX2TS U959 ( .A(\addr_calc/iir_read_calc/count[12] ), .Y(\add_x_22_4/n74 )
         );
  CLKBUFX2TS U960 ( .A(\addr_calc/iir_read_calc/count[10] ), .Y(n1909) );
  CLKBUFX2TS U961 ( .A(\addr_calc/fir_read_calc/count[1] ), .Y(n1910) );
  INVX2TS U962 ( .A(n1766), .Y(n1774) );
  INVX2TS U963 ( .A(n1765), .Y(n1769) );
  OAI2BB1X1TS U964 ( .A0N(n1533), .A1N(n1589), .B0(\add_x_19_5/n37 ), .Y(n1534) );
  NOR2BX1TS U965 ( .AN(n2629), .B(\add_x_19_5/n36 ), .Y(n1532) );
  INVX2TS U966 ( .A(n1765), .Y(n1768) );
  NOR2BX1TS U967 ( .AN(\add_x_19_4/n37 ), .B(\add_x_19_4/n36 ), .Y(n1640) );
  INVX2TS U968 ( .A(\add_x_19_4/n40 ), .Y(n1583) );
  OA21XLTS U969 ( .A0(\add_x_19_4/n36 ), .A1(n1583), .B0(\add_x_19_4/n37 ), 
        .Y(n1585) );
  NOR2BX1TS U970 ( .AN(n2634), .B(\add_x_19_4/n36 ), .Y(n1584) );
  INVX2TS U971 ( .A(\add_x_19_5/n42 ), .Y(n1589) );
  INVX2TS U972 ( .A(\add_x_19_2/n42 ), .Y(n1559) );
  INVX2TS U973 ( .A(n1766), .Y(n1773) );
  INVX2TS U974 ( .A(n1765), .Y(n1767) );
  NOR2X1TS U975 ( .A(n1297), .B(n1298), .Y(n2793) );
  INVX2TS U976 ( .A(n1820), .Y(n1827) );
  INVX2TS U977 ( .A(\addr_calc/fir_write_calc/count[18] ), .Y(n2005) );
  INVX2TS U978 ( .A(n1720), .Y(n1723) );
  INVX2TS U979 ( .A(\addr_calc/fir_read_calc/count[21] ), .Y(n1878) );
  BUFX8TS U980 ( .A(n2809), .Y(n1741) );
  INVX2TS U981 ( .A(n1820), .Y(n1824) );
  NOR2X1TS U982 ( .A(\addr_calc/iir_read_calc/count[5] ), .B(n2483), .Y(
        \add_x_19_4/n170 ) );
  NAND2X1TS U983 ( .A(n2426), .B(\addr_calc/iir_read_calc/count[14] ), .Y(
        \add_x_19_4/n124 ) );
  NAND2X1TS U984 ( .A(n1999), .B(n2408), .Y(\add_x_19_3/n132 ) );
  NOR2X1TS U985 ( .A(n1690), .B(n2424), .Y(\add_x_19_2/n123 ) );
  NAND2X1TS U986 ( .A(n2011), .B(n2462), .Y(\add_x_19_1/n67 ) );
  NOR2X1TS U987 ( .A(n2043), .B(n2426), .Y(\add_x_19_0/n123 ) );
  NAND2X1TS U988 ( .A(\addr_calc/iir_write_calc/count[16] ), .B(n2401), .Y(
        \add_x_19_5/n111 ) );
  NOR2X1TS U989 ( .A(n1992), .B(n2429), .Y(\add_x_19_3/n165 ) );
  NAND2X1TS U990 ( .A(n1995), .B(n2472), .Y(\add_x_19_3/n155 ) );
  NOR2X1TS U991 ( .A(\addr_calc/fft_write_calc/count[6] ), .B(n2428), .Y(
        \add_x_19_1/n165 ) );
  NOR2X2TS U992 ( .A(n1666), .B(n2422), .Y(\add_x_19_0/n162 ) );
  NOR2X1TS U993 ( .A(n1902), .B(n2436), .Y(\add_x_19_4/n181 ) );
  INVX2TS U994 ( .A(n2066), .Y(n2060) );
  INVX4TS U995 ( .A(\DP_OP_158_296_6262/n2060 ), .Y(\DP_OP_158_296_6262/n829 )
         );
  INVX2TS U996 ( .A(n2063), .Y(n1861) );
  INVX2TS U997 ( .A(n2584), .Y(n2588) );
  CLKBUFX2TS U998 ( .A(\addr_calc/fir_write_calc/count[25] ), .Y(n1894) );
  XOR2X1TS U999 ( .A(\DP_OP_158_296_6262/n2020 ), .B(n1680), .Y(n2596) );
  INVX6TS U1000 ( .A(\DP_OP_158_296_6262/n2054 ), .Y(n1718) );
  INVX6TS U1001 ( .A(\DP_OP_158_296_6262/n2056 ), .Y(\DP_OP_158_296_6262/n833 ) );
  INVX2TS U1002 ( .A(n1930), .Y(n1667) );
  CLKBUFX2TS U1003 ( .A(\addr_calc/fft_write_calc/count[14] ), .Y(n2021) );
  INVX2TS U1004 ( .A(n1497), .Y(\DP_OP_159_297_3515/n880 ) );
  NAND2BX1TS U1005 ( .AN(\add_x_19_2/n86 ), .B(\add_x_19_2/n87 ), .Y(n1569) );
  NAND2BX1TS U1006 ( .AN(\add_x_19_1/n36 ), .B(n1555), .Y(n1550) );
  AOI2BB2X1TS U1007 ( .B0(n1552), .B1(\add_x_19_1/n36 ), .A0N(\add_x_19_1/n37 ), .A1N(n1554), .Y(n1553) );
  XNOR2X1TS U1008 ( .A(\add_x_19_1/n88 ), .B(\add_x_19_1/n11 ), .Y(
        \addr_calc/fft_write_addr[21] ) );
  NAND2BX1TS U1009 ( .AN(n1543), .B(n1748), .Y(n1542) );
  NAND2BX1TS U1010 ( .AN(n1566), .B(n1772), .Y(n1565) );
  XNOR2X1TS U1011 ( .A(\add_x_22_5/n58 ), .B(\add_x_22_5/n57 ), .Y(n1566) );
  XNOR2X1TS U1012 ( .A(n1575), .B(n1948), .Y(n1574) );
  XNOR2X1TS U1013 ( .A(\add_x_22_3/n75 ), .B(n2000), .Y(n1647) );
  XNOR2X2TS U1014 ( .A(n1578), .B(\addr_calc/iir_read_calc/count[27] ), .Y(
        n1577) );
  NAND2BX1TS U1015 ( .AN(\add_x_19_2/n78 ), .B(\add_x_19_2/n79 ), .Y(n1597) );
  XNOR2X1TS U1016 ( .A(\add_x_22_3/n110 ), .B(\add_x_22_3/n109 ), .Y(n1616) );
  OAI2BB2X2TS U1017 ( .B0(n1740), .B1(\add_x_22_5/n80 ), .A0N(n1771), .A1N(
        \addr_calc/iir_write_calc/counter/N54 ), .Y(n991) );
  NAND2X1TS U1018 ( .A(n1752), .B(n1621), .Y(n1620) );
  XNOR2X1TS U1019 ( .A(n1622), .B(\add_x_22_0/n80 ), .Y(n1621) );
  XNOR2X1TS U1020 ( .A(\add_x_22_0/n102 ), .B(n1610), .Y(n1609) );
  XNOR2X1TS U1021 ( .A(\add_x_22_0/n110 ), .B(\add_x_22_0/n109 ), .Y(n1644) );
  XNOR2X1TS U1022 ( .A(\add_x_22_0/n58 ), .B(\add_x_22_0/n57 ), .Y(n1639) );
  XNOR2X1TS U1023 ( .A(\add_x_22_0/n50 ), .B(n2569), .Y(n1637) );
  XNOR2X1TS U1024 ( .A(\add_x_22_0/n16 ), .B(n2575), .Y(n1631) );
  XNOR2X1TS U1025 ( .A(\add_x_22_4/n16 ), .B(n1572), .Y(n1571) );
  OAI2BB1X1TS U1026 ( .A0N(n2582), .A1N(n1674), .B0(n1612), .Y(n1072) );
  XNOR2X1TS U1027 ( .A(\add_x_22_2/n16 ), .B(n1614), .Y(n1613) );
  INVX2TS U1028 ( .A(\add_x_22_2/n15 ), .Y(n1614) );
  NAND2BX1TS U1029 ( .AN(\add_x_19_5/n120 ), .B(\add_x_19_5/n121 ), .Y(n1537)
         );
  NOR2BX1TS U1030 ( .AN(\add_x_19_0/n37 ), .B(\add_x_19_0/n36 ), .Y(n1544) );
  NOR2BX1TS U1031 ( .AN(\add_x_19_3/n37 ), .B(\add_x_19_3/n36 ), .Y(n1538) );
  NAND2BX1TS U1032 ( .AN(\add_x_19_5/n58 ), .B(n1607), .Y(n1603) );
  XNOR2X1TS U1033 ( .A(\add_x_22_3/n41 ), .B(n2009), .Y(n1619) );
  NAND2X1TS U1034 ( .A(n1752), .B(n1628), .Y(n1627) );
  XNOR2X1TS U1035 ( .A(n1629), .B(n1953), .Y(n1628) );
  XNOR2X1TS U1036 ( .A(n1657), .B(n2043), .Y(\DP_OP_158_296_6262/n1149 ) );
  XNOR2X2TS U1037 ( .A(\DP_OP_158_296_6262/n838 ), .B(
        \addr_calc/fft_read_calc/count[21] ), .Y(\DP_OP_158_296_6262/n1055 )
         );
  XNOR2X1TS U1038 ( .A(n2594), .B(\addr_calc/fft_read_calc/count[16] ), .Y(
        \DP_OP_158_296_6262/n1124 ) );
  XNOR2X2TS U1039 ( .A(\DP_OP_159_297_3515/n885 ), .B(n2324), .Y(n2614) );
  XNOR2X2TS U1040 ( .A(\DP_OP_159_297_3515/n1044 ), .B(
        \DP_OP_159_297_3515/n876 ), .Y(n2622) );
  XNOR2X2TS U1041 ( .A(n2613), .B(n1839), .Y(n1624) );
  CLKBUFX2TS U1042 ( .A(n1518), .Y(n2344) );
  NOR2X1TS U1043 ( .A(\DP_OP_159_297_3515/n1012 ), .B(
        \DP_OP_159_297_3515/n991 ), .Y(\DP_OP_159_297_3515/n990 ) );
  NOR2X1TS U1044 ( .A(\DP_OP_158_296_6262/n2020 ), .B(n1680), .Y(
        \DP_OP_158_296_6262/n2015 ) );
  NAND2X1TS U1045 ( .A(n1783), .B(\DP_OP_158_296_6262/n1842 ), .Y(
        \DP_OP_158_296_6262/n1841 ) );
  NOR2X1TS U1046 ( .A(\DP_OP_158_296_6262/n1946 ), .B(n1831), .Y(
        \DP_OP_158_296_6262/n1938 ) );
  INVX2TS U1047 ( .A(n1508), .Y(n2343) );
  INVX2TS U1048 ( .A(n2342), .Y(n1464) );
  BUFX4TS U1049 ( .A(n1482), .Y(n1831) );
  INVX4TS U1050 ( .A(\DP_OP_159_297_3515/n1133 ), .Y(\DP_OP_159_297_3515/n792 ) );
  OAI21XLTS U1051 ( .A0(\add_x_19_5/n120 ), .A1(\add_x_19_5/n124 ), .B0(
        \add_x_19_5/n121 ), .Y(n1271) );
  AOI21X1TS U1052 ( .A0(\add_x_19_5/n127 ), .A1(\add_x_19_5/n118 ), .B0(n1271), 
        .Y(\add_x_19_5/n117 ) );
  OAI21X1TS U1053 ( .A0(\add_x_19_1/n139 ), .A1(\add_x_19_1/n145 ), .B0(
        \add_x_19_1/n140 ), .Y(n1272) );
  AOI21X1TS U1054 ( .A0(\add_x_19_1/n150 ), .A1(\add_x_19_1/n137 ), .B0(n1272), 
        .Y(\add_x_19_1/n136 ) );
  NOR2X1TS U1055 ( .A(\add_x_22_3/n94 ), .B(n1273), .Y(\add_x_22_3/n59 ) );
  NAND4BX1TS U1056 ( .AN(\add_x_22_0/n69 ), .B(n2043), .C(n1689), .D(
        \add_x_22_0/n77 ), .Y(n1274) );
  NOR2X1TS U1057 ( .A(\add_x_22_0/n94 ), .B(n1274), .Y(\add_x_22_0/n59 ) );
  NAND3X1TS U1058 ( .A(\addr_calc/iir_read_calc/count[15] ), .B(
        \addr_calc/iir_read_calc/count[14] ), .C(\add_x_22_4/n77 ), .Y(n1275)
         );
  NOR3X1TS U1059 ( .A(\add_x_22_4/n94 ), .B(\add_x_22_4/n69 ), .C(n1275), .Y(
        \add_x_22_4/n59 ) );
  NAND3X1TS U1060 ( .A(n1890), .B(n1690), .C(\add_x_22_2/n77 ), .Y(n1276) );
  NOR3X1TS U1061 ( .A(\add_x_22_2/n94 ), .B(\add_x_22_2/n69 ), .C(n1276), .Y(
        \add_x_22_2/n59 ) );
  NAND2BX1TS U1062 ( .AN(\add_x_19_2/n36 ), .B(\add_x_19_2/n37 ), .Y(n1277) );
  XOR2X2TS U1063 ( .A(\add_x_19_2/n38 ), .B(n1277), .Y(
        \addr_calc/fir_read_addr[30] ) );
  NAND2BX1TS U1064 ( .AN(\add_x_19_0/n66 ), .B(\add_x_19_0/n67 ), .Y(n1278) );
  XOR2X1TS U1065 ( .A(\add_x_19_0/n68 ), .B(n1278), .Y(
        \addr_calc/fft_read_addr[24] ) );
  NAND2BX1TS U1066 ( .AN(\add_x_19_4/n89 ), .B(\add_x_19_4/n90 ), .Y(n1279) );
  XOR2X1TS U1067 ( .A(\add_x_19_4/n91 ), .B(n1279), .Y(
        \addr_calc/iir_read_addr[20] ) );
  NAND2BX1TS U1068 ( .AN(\add_x_19_2/n165 ), .B(\add_x_19_2/n166 ), .Y(n1280)
         );
  XOR2X1TS U1069 ( .A(\add_x_19_2/n167 ), .B(n1280), .Y(
        \addr_calc/fir_read_addr[6] ) );
  NAND2BX1TS U1070 ( .AN(\add_x_19_1/n165 ), .B(\add_x_19_1/n166 ), .Y(n1281)
         );
  XOR2X1TS U1071 ( .A(\add_x_19_1/n167 ), .B(n1281), .Y(
        \addr_calc/fft_write_addr[6] ) );
  OAI21XLTS U1072 ( .A0(\add_x_19_3/n154 ), .A1(\add_x_19_3/n156 ), .B0(
        \add_x_19_3/n155 ), .Y(n1282) );
  CLKINVX1TS U1073 ( .A(\add_x_19_3/n152 ), .Y(n1283) );
  OAI21XLTS U1074 ( .A0(\add_x_19_3/n151 ), .A1(n1283), .B0(n1282), .Y(n1284)
         );
  OAI31XLTS U1075 ( .A0(\add_x_19_3/n151 ), .A1(n1282), .A2(n1283), .B0(n1284), 
        .Y(\addr_calc/fir_write_addr[9] ) );
  OAI21X1TS U1076 ( .A0(\add_x_19_4/n184 ), .A1(\add_x_19_4/n186 ), .B0(
        \add_x_19_4/n185 ), .Y(n1285) );
  CLKINVX1TS U1077 ( .A(\add_x_19_4/n182 ), .Y(n1286) );
  OAI21X1TS U1078 ( .A0(\add_x_19_4/n181 ), .A1(n1286), .B0(n1285), .Y(n1287)
         );
  OAI31X1TS U1079 ( .A0(\add_x_19_4/n181 ), .A1(n1285), .A2(n1286), .B0(n1287), 
        .Y(\addr_calc/iir_read_addr[3] ) );
  OA21XLTS U1080 ( .A0(n2578), .A1(n2394), .B0(\add_x_19_5/n191 ), .Y(
        \addr_calc/iir_write_addr[0] ) );
  NAND2BX1TS U1081 ( .AN(\add_x_22_3/n26 ), .B(\add_x_22_3/n59 ), .Y(
        \add_x_22_3/n24 ) );
  NAND3X1TS U1082 ( .A(\addr_calc/iir_write_calc/count[15] ), .B(
        \addr_calc/iir_write_calc/count[14] ), .C(\add_x_22_5/n77 ), .Y(n1288)
         );
  NOR3X1TS U1083 ( .A(\add_x_22_5/n94 ), .B(\add_x_22_5/n69 ), .C(n1288), .Y(
        \add_x_22_5/n59 ) );
  NOR4XLTS U1084 ( .A(n2022), .B(n1927), .C(n1976), .D(
        \addr_calc/fft_write_calc/count[16] ), .Y(n1289) );
  NOR4XLTS U1085 ( .A(n2023), .B(n2035), .C(
        \addr_calc/fft_write_calc/count[11] ), .D(n1932), .Y(n1290) );
  NAND4X1TS U1086 ( .A(n1289), .B(n1290), .C(n847), .D(n846), .Y(n1291) );
  NAND4X1TS U1087 ( .A(n845), .B(n844), .C(n843), .D(n842), .Y(n1292) );
  NOR2X1TS U1088 ( .A(n1291), .B(n1292), .Y(n2796) );
  CLKINVX1TS U1089 ( .A(n1607), .Y(n1293) );
  CLKINVX1TS U1090 ( .A(n1473), .Y(n1294) );
  AOI32X1TS U1091 ( .A0(\add_x_19_5/n58 ), .A1(n1293), .A2(\add_x_19_5/n59 ), 
        .B0(n1607), .B1(n1294), .Y(n1606) );
  NOR4XLTS U1092 ( .A(n1970), .B(\addr_calc/fft_read_calc/count[12] ), .C(
        n2058), .D(n1972), .Y(n1295) );
  NOR4XLTS U1093 ( .A(\addr_calc/fft_read_calc/count[15] ), .B(
        \addr_calc/fft_read_calc/count[14] ), .C(n1967), .D(n2554), .Y(n1296)
         );
  NAND4X1TS U1094 ( .A(n832), .B(n833), .C(n1295), .D(n1296), .Y(n1297) );
  NAND4X1TS U1095 ( .A(n828), .B(n829), .C(n830), .D(n831), .Y(n1298) );
  AOI21X1TS U1096 ( .A0(\add_x_19_3/n73 ), .A1(\add_x_19_3/n46 ), .B0(
        \add_x_19_3/n47 ), .Y(n1299) );
  OAI2BB1X2TS U1097 ( .A0N(n1470), .A1N(n1676), .B0(n1299), .Y(
        \add_x_19_3/n43 ) );
  OAI21X1TS U1098 ( .A0(\add_x_19_3/n131 ), .A1(\add_x_19_3/n133 ), .B0(
        \add_x_19_3/n132 ), .Y(n1300) );
  CLKINVX1TS U1099 ( .A(\add_x_19_3/n129 ), .Y(n1301) );
  OAI21XLTS U1100 ( .A0(\add_x_19_3/n128 ), .A1(n1301), .B0(n1300), .Y(n1302)
         );
  OAI2BB1X1TS U1101 ( .A0N(n1818), .A1N(\add_x_19_5/n219 ), .B0(
        \add_x_19_5/n176 ), .Y(n1303) );
  CLKINVX1TS U1102 ( .A(\add_x_19_5/n171 ), .Y(n1304) );
  OAI21XLTS U1103 ( .A0(\add_x_19_5/n170 ), .A1(n1304), .B0(n1303), .Y(n1305)
         );
  OAI31XLTS U1104 ( .A0(\add_x_19_5/n170 ), .A1(n1303), .A2(n1304), .B0(n1305), 
        .Y(\addr_calc/iir_write_addr[5] ) );
  OAI2BB1X2TS U1105 ( .A0N(\add_x_19_5/n146 ), .A1N(\add_x_19_5/n213 ), .B0(
        \add_x_19_5/n145 ), .Y(n1306) );
  CLKINVX1TS U1106 ( .A(\add_x_19_5/n140 ), .Y(n1307) );
  OAI21X1TS U1107 ( .A0(\add_x_19_5/n139 ), .A1(n1307), .B0(n1306), .Y(n1308)
         );
  OAI31X1TS U1108 ( .A0(\add_x_19_5/n139 ), .A1(n1306), .A2(n1307), .B0(n1308), 
        .Y(\addr_calc/iir_write_addr[11] ) );
  NAND2BX1TS U1109 ( .AN(\add_x_19_5/n66 ), .B(\add_x_19_5/n67 ), .Y(n1309) );
  XOR2X1TS U1110 ( .A(\add_x_19_5/n68 ), .B(n1309), .Y(
        \addr_calc/iir_write_addr[24] ) );
  NAND2BX1TS U1111 ( .AN(\add_x_19_0/n165 ), .B(\add_x_19_0/n166 ), .Y(n1310)
         );
  XOR2X1TS U1112 ( .A(\add_x_19_0/n167 ), .B(n1310), .Y(
        \addr_calc/fft_read_addr[6] ) );
  OAI2BB1X1TS U1113 ( .A0N(\add_x_19_0/n146 ), .A1N(\add_x_19_0/n213 ), .B0(
        \add_x_19_0/n145 ), .Y(n1311) );
  CLKINVX1TS U1114 ( .A(\add_x_19_0/n140 ), .Y(n1312) );
  OAI21X1TS U1115 ( .A0(\add_x_19_0/n139 ), .A1(n1312), .B0(n1311), .Y(n1313)
         );
  OAI31X1TS U1116 ( .A0(\add_x_19_0/n139 ), .A1(n1311), .A2(n1312), .B0(n1313), 
        .Y(\addr_calc/fft_read_addr[11] ) );
  OAI21XLTS U1117 ( .A0(\add_x_19_3/n184 ), .A1(\add_x_19_3/n186 ), .B0(
        \add_x_19_3/n185 ), .Y(n1314) );
  CLKINVX1TS U1118 ( .A(\add_x_19_3/n182 ), .Y(n1315) );
  OAI21X1TS U1119 ( .A0(\add_x_19_3/n181 ), .A1(n1315), .B0(n1314), .Y(n1316)
         );
  OAI31X1TS U1120 ( .A0(\add_x_19_3/n181 ), .A1(n1314), .A2(n1315), .B0(n1316), 
        .Y(\addr_calc/fir_write_addr[3] ) );
  OA21XLTS U1121 ( .A0(n2580), .A1(n2393), .B0(\add_x_19_4/n191 ), .Y(
        \addr_calc/iir_read_addr[0] ) );
  NOR4XLTS U1122 ( .A(n2107), .B(n2088), .C(n2080), .D(n1803), .Y(n1317) );
  NOR4XLTS U1123 ( .A(n2112), .B(n2097), .C(n2082), .D(n2101), .Y(n1318) );
  NOR4BBX1TS U1124 ( .AN(n2108), .BN(n2093), .C(n2078), .D(n2099), .Y(n1319)
         );
  NAND4X1TS U1125 ( .A(n1317), .B(n802), .C(n1318), .D(n1319), .Y(n908) );
  NAND4BX1TS U1126 ( .AN(\add_x_22_5/n103 ), .B(\add_x_22_5/n111 ), .C(n1683), 
        .D(\addr_calc/iir_write_calc/count[6] ), .Y(\add_x_22_5/n94 ) );
  NAND4BX1TS U1127 ( .AN(\add_x_22_3/n103 ), .B(\add_x_22_3/n111 ), .C(n1869), 
        .D(n1993), .Y(\add_x_22_3/n94 ) );
  NAND2BX1TS U1128 ( .AN(\add_x_22_2/n26 ), .B(\add_x_22_2/n59 ), .Y(
        \add_x_22_2/n24 ) );
  NAND2BX1TS U1129 ( .AN(\add_x_22_4/n87 ), .B(\add_x_22_4/n93 ), .Y(
        \add_x_22_4/n85 ) );
  CLKINVX1TS U1130 ( .A(n1640), .Y(n1320) );
  OAI32X1TS U1131 ( .A0(n1320), .A1(\add_x_19_4/n40 ), .A2(n2634), .B0(n1640), 
        .B1(n1583), .Y(n1582) );
  NAND2BX1TS U1132 ( .AN(\add_x_19_1/n58 ), .B(\add_x_19_1/n59 ), .Y(n1321) );
  NAND2BX1TS U1133 ( .AN(\add_x_19_1/n100 ), .B(\add_x_19_1/n101 ), .Y(n1322)
         );
  XOR2X1TS U1134 ( .A(\add_x_19_1/n102 ), .B(n1322), .Y(
        \addr_calc/fft_write_addr[18] ) );
  NAND2BX1TS U1135 ( .AN(\add_x_19_5/n81 ), .B(\add_x_19_5/n82 ), .Y(n1323) );
  XOR2X1TS U1136 ( .A(\add_x_19_5/n83 ), .B(n1323), .Y(
        \addr_calc/iir_write_addr[22] ) );
  XNOR2X1TS U1137 ( .A(\add_x_22_1/n117 ), .B(\add_x_22_1/n118 ), .Y(n1324) );
  AO22X4TS U1138 ( .A0(n2662), .A1(n2032), .B0(n1724), .B1(n1324), .Y(n1064)
         );
  NAND2BX1TS U1139 ( .AN(\add_x_19_2/n58 ), .B(\add_x_19_2/n59 ), .Y(n1325) );
  NAND2BX1TS U1140 ( .AN(\add_x_19_5/n154 ), .B(\add_x_19_5/n155 ), .Y(n1326)
         );
  XOR2X1TS U1141 ( .A(\add_x_19_5/n156 ), .B(n1326), .Y(
        \addr_calc/iir_write_addr[8] ) );
  NAND2BX1TS U1142 ( .AN(\add_x_19_5/n131 ), .B(\add_x_19_5/n132 ), .Y(n1327)
         );
  XOR2X1TS U1143 ( .A(\add_x_19_5/n133 ), .B(n1327), .Y(
        \addr_calc/iir_write_addr[12] ) );
  OAI2BB1X1TS U1144 ( .A0N(\add_x_19_3/n146 ), .A1N(\add_x_19_3/n213 ), .B0(
        \add_x_19_3/n145 ), .Y(n1328) );
  CLKINVX1TS U1145 ( .A(\add_x_19_3/n140 ), .Y(n1329) );
  OAI21X1TS U1146 ( .A0(\add_x_19_3/n139 ), .A1(n1329), .B0(n1328), .Y(n1330)
         );
  OAI31XLTS U1147 ( .A0(\add_x_19_3/n139 ), .A1(n1328), .A2(n1329), .B0(n1330), 
        .Y(\addr_calc/fir_write_addr[11] ) );
  OAI2BB1X2TS U1148 ( .A0N(n1676), .A1N(\add_x_19_3/n207 ), .B0(
        \add_x_19_3/n111 ), .Y(n1331) );
  CLKINVX1TS U1149 ( .A(\add_x_19_3/n106 ), .Y(n1332) );
  OAI21X1TS U1150 ( .A0(\add_x_19_3/n105 ), .A1(n1332), .B0(n1331), .Y(n1333)
         );
  OAI31X1TS U1151 ( .A0(\add_x_19_3/n105 ), .A1(n1331), .A2(n1332), .B0(n1333), 
        .Y(\addr_calc/fir_write_addr[17] ) );
  NAND2BX1TS U1152 ( .AN(\add_x_19_3/n66 ), .B(\add_x_19_3/n67 ), .Y(n1334) );
  XOR2X1TS U1153 ( .A(\add_x_19_3/n68 ), .B(n1334), .Y(
        \addr_calc/fir_write_addr[24] ) );
  OAI2BB1X1TS U1154 ( .A0N(\add_x_19_2/n177 ), .A1N(\add_x_19_2/n219 ), .B0(
        \add_x_19_2/n176 ), .Y(n1335) );
  CLKINVX1TS U1155 ( .A(\add_x_19_2/n171 ), .Y(n1336) );
  OAI21XLTS U1156 ( .A0(\add_x_19_2/n170 ), .A1(n1336), .B0(n1335), .Y(n1337)
         );
  OAI31XLTS U1157 ( .A0(\add_x_19_2/n170 ), .A1(n1335), .A2(n1336), .B0(n1337), 
        .Y(\addr_calc/fir_read_addr[5] ) );
  OAI21X1TS U1158 ( .A0(\add_x_19_4/n165 ), .A1(\add_x_19_4/n167 ), .B0(
        \add_x_19_4/n166 ), .Y(n1338) );
  CLKINVX1TS U1159 ( .A(\add_x_19_4/n163 ), .Y(n1339) );
  OAI21X1TS U1160 ( .A0(\add_x_19_4/n162 ), .A1(n1339), .B0(n1338), .Y(n1340)
         );
  OAI31X1TS U1161 ( .A0(\add_x_19_4/n162 ), .A1(n1338), .A2(n1339), .B0(n1340), 
        .Y(\addr_calc/iir_read_addr[7] ) );
  OAI21X1TS U1162 ( .A0(\add_x_19_2/n154 ), .A1(\add_x_19_2/n156 ), .B0(
        \add_x_19_2/n155 ), .Y(n1341) );
  INVXLTS U1163 ( .A(\add_x_19_2/n152 ), .Y(n1342) );
  OAI21XLTS U1164 ( .A0(\add_x_19_2/n151 ), .A1(n1342), .B0(n1341), .Y(n1343)
         );
  OAI31XLTS U1165 ( .A0(\add_x_19_2/n151 ), .A1(n1341), .A2(n1342), .B0(n1343), 
        .Y(\addr_calc/fir_read_addr[9] ) );
  NAND2BX1TS U1166 ( .AN(\add_x_19_5/n184 ), .B(\add_x_19_5/n185 ), .Y(n1344)
         );
  XOR2X1TS U1167 ( .A(\add_x_19_5/n186 ), .B(n1344), .Y(
        \addr_calc/iir_write_addr[2] ) );
  NAND2BX1TS U1168 ( .AN(\add_x_19_2/n188 ), .B(\add_x_19_2/n189 ), .Y(n1345)
         );
  XOR2X1TS U1169 ( .A(\add_x_19_2/n191 ), .B(n1345), .Y(
        \addr_calc/fir_read_addr[1] ) );
  OAI21X1TS U1170 ( .A0(\add_x_19_2/n184 ), .A1(\add_x_19_2/n186 ), .B0(
        \add_x_19_2/n185 ), .Y(n1346) );
  CLKINVX1TS U1171 ( .A(\add_x_19_2/n182 ), .Y(n1347) );
  OAI21X1TS U1172 ( .A0(\add_x_19_2/n181 ), .A1(n1347), .B0(n1346), .Y(n1348)
         );
  OAI31X1TS U1173 ( .A0(\add_x_19_2/n181 ), .A1(n1346), .A2(n1347), .B0(n1348), 
        .Y(\addr_calc/fir_read_addr[3] ) );
  OA21XLTS U1174 ( .A0(n1986), .A1(n2394), .B0(\add_x_19_3/n191 ), .Y(
        \addr_calc/fir_write_addr[0] ) );
  NAND4BX1TS U1175 ( .AN(\add_x_22_1/n69 ), .B(n2021), .C(
        \addr_calc/fft_write_calc/count[15] ), .D(\add_x_22_1/n77 ), .Y(n1349)
         );
  NOR2X2TS U1176 ( .A(\add_x_22_1/n94 ), .B(n1349), .Y(\add_x_22_1/n59 ) );
  NAND2BX1TS U1177 ( .AN(\add_x_22_5/n26 ), .B(\add_x_22_5/n59 ), .Y(
        \add_x_22_5/n24 ) );
  NAND4BX1TS U1178 ( .AN(\add_x_22_4/n103 ), .B(\add_x_22_4/n111 ), .C(n1905), 
        .D(\addr_calc/iir_read_calc/count[6] ), .Y(\add_x_22_4/n94 ) );
  NAND2BX1TS U1179 ( .AN(\add_x_22_0/n87 ), .B(\add_x_22_0/n93 ), .Y(
        \add_x_22_0/n85 ) );
  AND4X1TS U1180 ( .A(n1799), .B(n1805), .C(instruction[29]), .D(
        instruction[30]), .Y(n1350) );
  AND3X1TS U1181 ( .A(instruction[31]), .B(n1801), .C(n1350), .Y(n802) );
  NAND2BX1TS U1182 ( .AN(\add_x_19_0/n100 ), .B(\add_x_19_0/n101 ), .Y(n1351)
         );
  XOR2X1TS U1183 ( .A(\add_x_19_0/n102 ), .B(n1351), .Y(
        \addr_calc/fft_read_addr[18] ) );
  NAND2BX1TS U1184 ( .AN(\add_x_19_2/n81 ), .B(\add_x_19_2/n82 ), .Y(n1352) );
  XOR2X1TS U1185 ( .A(\add_x_19_2/n83 ), .B(n1352), .Y(
        \addr_calc/fir_read_addr[22] ) );
  XNOR2X1TS U1186 ( .A(\addr_calc/fft_write_calc/count[0] ), .B(
        \add_x_22_1/n121 ), .Y(n1353) );
  AO22X4TS U1187 ( .A0(n2662), .A1(n1941), .B0(n1721), .B1(n1353), .Y(n1065)
         );
  NAND2BX1TS U1188 ( .AN(\add_x_19_5/n58 ), .B(n1473), .Y(n1354) );
  XOR2X1TS U1189 ( .A(\add_x_19_5/n60 ), .B(n1354), .Y(
        \addr_calc/iir_write_addr[26] ) );
  NAND2BX1TS U1190 ( .AN(\add_x_19_4/n58 ), .B(\add_x_19_4/n59 ), .Y(n1355) );
  XOR2X2TS U1191 ( .A(\add_x_19_4/n60 ), .B(n1355), .Y(
        \addr_calc/iir_read_addr[26] ) );
  OAI2BB1X4TS U1192 ( .A0N(n1584), .A1N(\add_x_19_4/n43 ), .B0(n1585), .Y(
        n1356) );
  OAI2BB1X1TS U1193 ( .A0N(\addr_calc/iir_read_calc/count[31] ), .A1N(n2381), 
        .B0(n1586), .Y(n1357) );
  AOI21X1TS U1194 ( .A0(\add_x_19_5/n43 ), .A1(n2629), .B0(n1589), .Y(n1358)
         );
  NAND2X1TS U1195 ( .A(n1533), .B(\add_x_19_5/n37 ), .Y(n1359) );
  XOR2X1TS U1196 ( .A(n1358), .B(n1359), .Y(\addr_calc/iir_write_addr[30] ) );
  NAND2BX1TS U1197 ( .AN(\add_x_19_5/n123 ), .B(\add_x_19_5/n124 ), .Y(n1360)
         );
  XOR2X1TS U1198 ( .A(\add_x_19_5/n125 ), .B(n1360), .Y(
        \addr_calc/iir_write_addr[14] ) );
  NAND2BX1TS U1199 ( .AN(\add_x_19_5/n89 ), .B(\add_x_19_5/n90 ), .Y(n1361) );
  XOR2X1TS U1200 ( .A(\add_x_19_5/n91 ), .B(n1361), .Y(
        \addr_calc/iir_write_addr[20] ) );
  NAND2BX1TS U1201 ( .AN(\add_x_19_4/n154 ), .B(\add_x_19_4/n155 ), .Y(n1362)
         );
  XOR2X1TS U1202 ( .A(\add_x_19_4/n156 ), .B(n1362), .Y(
        \addr_calc/iir_read_addr[8] ) );
  NAND2BX1TS U1203 ( .AN(\add_x_19_2/n131 ), .B(\add_x_19_2/n132 ), .Y(n1363)
         );
  XOR2X1TS U1204 ( .A(\add_x_19_2/n133 ), .B(n1363), .Y(
        \addr_calc/fir_read_addr[12] ) );
  NAND2BX1TS U1205 ( .AN(\add_x_19_2/n66 ), .B(\add_x_19_2/n67 ), .Y(n1364) );
  XOR2X1TS U1206 ( .A(\add_x_19_2/n68 ), .B(n1364), .Y(
        \addr_calc/fir_read_addr[24] ) );
  NAND2BX1TS U1207 ( .AN(\add_x_19_0/n184 ), .B(\add_x_19_0/n185 ), .Y(n1365)
         );
  XOR2X1TS U1208 ( .A(\add_x_19_0/n186 ), .B(n1365), .Y(
        \addr_calc/fft_read_addr[2] ) );
  CLKINVX1TS U1209 ( .A(\add_x_19_0/n171 ), .Y(n1366) );
  OAI2BB1X1TS U1210 ( .A0N(\add_x_19_0/n177 ), .A1N(\add_x_19_0/n219 ), .B0(
        \add_x_19_0/n176 ), .Y(n1367) );
  OAI21XLTS U1211 ( .A0(\add_x_19_0/n170 ), .A1(n1366), .B0(n1367), .Y(n1368)
         );
  OAI31XLTS U1212 ( .A0(\add_x_19_0/n170 ), .A1(n1367), .A2(n1366), .B0(n1368), 
        .Y(\addr_calc/fft_read_addr[5] ) );
  OAI21X1TS U1213 ( .A0(\add_x_19_5/n165 ), .A1(\add_x_19_5/n167 ), .B0(
        \add_x_19_5/n166 ), .Y(n1369) );
  CLKINVX1TS U1214 ( .A(\add_x_19_5/n163 ), .Y(n1370) );
  OAI21XLTS U1215 ( .A0(\add_x_19_5/n162 ), .A1(n1370), .B0(n1369), .Y(n1371)
         );
  OAI31XLTS U1216 ( .A0(\add_x_19_5/n162 ), .A1(n1369), .A2(n1370), .B0(n1371), 
        .Y(\addr_calc/iir_write_addr[7] ) );
  NAND2X1TS U1217 ( .A(\add_x_19_3/n207 ), .B(\add_x_19_3/n111 ), .Y(n1372) );
  XNOR2X1TS U1218 ( .A(n1372), .B(n1676), .Y(\addr_calc/fir_write_addr[16] )
         );
  OAI21XLTS U1219 ( .A0(\add_x_19_1/n165 ), .A1(\add_x_19_1/n167 ), .B0(
        \add_x_19_1/n166 ), .Y(n1373) );
  CLKINVX1TS U1220 ( .A(\add_x_19_1/n163 ), .Y(n1374) );
  OAI21X1TS U1221 ( .A0(\add_x_19_1/n162 ), .A1(n1374), .B0(n1373), .Y(n1375)
         );
  OAI31X1TS U1222 ( .A0(\add_x_19_1/n162 ), .A1(n1373), .A2(n1374), .B0(n1375), 
        .Y(\addr_calc/fft_write_addr[7] ) );
  OAI21XLTS U1223 ( .A0(\add_x_19_1/n154 ), .A1(\add_x_19_1/n156 ), .B0(
        \add_x_19_1/n155 ), .Y(n1376) );
  CLKINVX1TS U1224 ( .A(\add_x_19_1/n152 ), .Y(n1377) );
  OAI21XLTS U1225 ( .A0(\add_x_19_1/n151 ), .A1(n1377), .B0(n1376), .Y(n1378)
         );
  OAI31X1TS U1226 ( .A0(\add_x_19_1/n151 ), .A1(n1376), .A2(n1377), .B0(n1378), 
        .Y(\addr_calc/fft_write_addr[9] ) );
  NAND2BX1TS U1227 ( .AN(\add_x_19_3/n188 ), .B(\add_x_19_3/n189 ), .Y(n1379)
         );
  XOR2X1TS U1228 ( .A(\add_x_19_3/n191 ), .B(n1379), .Y(
        \addr_calc/fir_write_addr[1] ) );
  OAI21X1TS U1229 ( .A0(\add_x_19_1/n184 ), .A1(\add_x_19_1/n186 ), .B0(
        \add_x_19_1/n185 ), .Y(n1380) );
  CLKINVX1TS U1230 ( .A(\add_x_19_1/n182 ), .Y(n1381) );
  OAI21XLTS U1231 ( .A0(\add_x_19_1/n181 ), .A1(n1381), .B0(n1380), .Y(n1382)
         );
  OAI31X1TS U1232 ( .A0(\add_x_19_1/n181 ), .A1(n1380), .A2(n1381), .B0(n1382), 
        .Y(\addr_calc/fft_write_addr[3] ) );
  OA21XLTS U1233 ( .A0(n2007), .A1(n2394), .B0(\add_x_19_2/n191 ), .Y(
        \addr_calc/fir_read_addr[0] ) );
  NAND4BX1TS U1234 ( .AN(\add_x_22_2/n35 ), .B(n2558), .C(n1691), .D(
        \add_x_22_2/n43 ), .Y(\add_x_22_2/n26 ) );
  NAND4BX1TS U1235 ( .AN(\add_x_22_0/n35 ), .B(
        \addr_calc/fft_read_calc/count[23] ), .C(
        \addr_calc/fft_read_calc/count[22] ), .D(\add_x_22_0/n43 ), .Y(
        \add_x_22_0/n26 ) );
  NAND2BX1TS U1236 ( .AN(\add_x_22_4/n26 ), .B(\add_x_22_4/n59 ), .Y(
        \add_x_22_4/n24 ) );
  NAND2BX1TS U1237 ( .AN(\add_x_22_1/n26 ), .B(\add_x_22_1/n59 ), .Y(
        \add_x_22_1/n24 ) );
  NAND2BX1TS U1238 ( .AN(\add_x_22_3/n87 ), .B(\add_x_22_3/n93 ), .Y(
        \add_x_22_3/n85 ) );
  NAND2BX1TS U1239 ( .AN(\add_x_22_2/n87 ), .B(\add_x_22_2/n93 ), .Y(
        \add_x_22_2/n85 ) );
  NAND2BX1TS U1240 ( .AN(n2311), .B(n902), .Y(n884) );
  XOR2X1TS U1241 ( .A(\add_x_22_4/n34 ), .B(n2031), .Y(n1383) );
  AO22X4TS U1242 ( .A0(n1708), .A1(n1383), .B0(n2031), .B1(n2651), .Y(n949) );
  AOI21X1TS U1243 ( .A0(\add_x_19_1/n207 ), .A1(\add_x_19_1/n112 ), .B0(
        \add_x_19_1/n109 ), .Y(n1384) );
  NAND2BX1TS U1244 ( .AN(\add_x_19_1/n105 ), .B(\add_x_19_1/n106 ), .Y(n1385)
         );
  XOR2X1TS U1245 ( .A(n1384), .B(n1385), .Y(\addr_calc/fft_write_addr[17] ) );
  NAND2BX1TS U1246 ( .AN(\add_x_19_1/n123 ), .B(\add_x_19_1/n124 ), .Y(n1386)
         );
  XOR2X1TS U1247 ( .A(\add_x_19_1/n125 ), .B(n1386), .Y(
        \addr_calc/fft_write_addr[14] ) );
  NAND2BX1TS U1248 ( .AN(\add_x_19_5/n100 ), .B(\add_x_19_5/n101 ), .Y(n1387)
         );
  XOR2X1TS U1249 ( .A(\add_x_19_5/n102 ), .B(n1387), .Y(
        \addr_calc/iir_write_addr[18] ) );
  NAND2BX1TS U1250 ( .AN(\add_x_19_4/n100 ), .B(\add_x_19_4/n101 ), .Y(n1388)
         );
  XOR2X1TS U1251 ( .A(\add_x_19_4/n102 ), .B(n1388), .Y(
        \addr_calc/iir_read_addr[18] ) );
  NOR2X1TS U1252 ( .A(\add_x_22_1/n84 ), .B(\add_x_22_1/n85 ), .Y(n1389) );
  XNOR2X1TS U1253 ( .A(n1389), .B(n1930), .Y(n1390) );
  AO22X4TS U1254 ( .A0(n2665), .A1(n1667), .B0(n1694), .B1(n1390), .Y(n1055)
         );
  NAND2BX1TS U1255 ( .AN(\add_x_19_3/n81 ), .B(\add_x_19_3/n82 ), .Y(n1391) );
  XOR2X1TS U1256 ( .A(\add_x_19_3/n83 ), .B(n1391), .Y(
        \addr_calc/fir_write_addr[22] ) );
  NAND2BX1TS U1257 ( .AN(\add_x_19_0/n58 ), .B(\add_x_19_0/n59 ), .Y(n1392) );
  XOR2X1TS U1258 ( .A(\add_x_19_0/n60 ), .B(n1392), .Y(
        \addr_calc/fft_read_addr[26] ) );
  NAND2BX1TS U1259 ( .AN(\add_x_19_0/n89 ), .B(\add_x_19_0/n90 ), .Y(n1393) );
  OAI2BB2X1TS U1260 ( .B0(n1476), .B1(n1394), .A0N(
        \addr_calc/fft_read_calc/count[0] ), .A1N(n1477), .Y(n1034) );
  NAND2X1TS U1261 ( .A(\add_x_22_3/n41 ), .B(n1669), .Y(n1395) );
  XOR2X1TS U1262 ( .A(n1891), .B(n1395), .Y(n1396) );
  AO22X4TS U1263 ( .A0(\addr_calc/fir_write_calc/count[21] ), .A1(n1260), .B0(
        n1762), .B1(n1396), .Y(n1109) );
  OAI2BB1X1TS U1264 ( .A0N(\add_x_19_4/n177 ), .A1N(\add_x_19_4/n219 ), .B0(
        \add_x_19_4/n176 ), .Y(n1397) );
  CLKINVX1TS U1265 ( .A(\add_x_19_4/n171 ), .Y(n1398) );
  OAI21X1TS U1266 ( .A0(\add_x_19_4/n170 ), .A1(n1398), .B0(n1397), .Y(n1399)
         );
  OAI31X1TS U1267 ( .A0(\add_x_19_4/n170 ), .A1(n1397), .A2(n1398), .B0(n1399), 
        .Y(\addr_calc/iir_read_addr[5] ) );
  NAND2BX1TS U1268 ( .AN(\add_x_19_4/n123 ), .B(\add_x_19_4/n124 ), .Y(n1400)
         );
  XOR2X1TS U1269 ( .A(\add_x_19_4/n125 ), .B(n1400), .Y(
        \addr_calc/iir_read_addr[14] ) );
  NAND2BX1TS U1270 ( .AN(\add_x_19_3/n131 ), .B(\add_x_19_3/n132 ), .Y(n1401)
         );
  XOR2X1TS U1271 ( .A(\add_x_19_3/n133 ), .B(n1401), .Y(
        \addr_calc/fir_write_addr[12] ) );
  AOI21X1TS U1272 ( .A0(\add_x_19_2/n146 ), .A1(\add_x_19_2/n213 ), .B0(
        \add_x_19_2/n143 ), .Y(n1402) );
  NAND2X1TS U1273 ( .A(\add_x_19_2/n212 ), .B(\add_x_19_2/n140 ), .Y(n1403) );
  XOR2X2TS U1274 ( .A(n1402), .B(n1403), .Y(\addr_calc/fir_read_addr[11] ) );
  NAND2BX1TS U1275 ( .AN(\add_x_19_2/n89 ), .B(\add_x_19_2/n90 ), .Y(n1404) );
  NAND2BX1TS U1276 ( .AN(\add_x_19_1/n154 ), .B(\add_x_19_1/n155 ), .Y(n1405)
         );
  NAND2BX1TS U1277 ( .AN(\add_x_19_1/n66 ), .B(\add_x_19_1/n67 ), .Y(n1406) );
  NAND2BX1TS U1278 ( .AN(\add_x_19_0/n131 ), .B(\add_x_19_0/n132 ), .Y(n1407)
         );
  XOR2X1TS U1279 ( .A(\add_x_19_0/n133 ), .B(n1407), .Y(
        \addr_calc/fft_read_addr[12] ) );
  NAND2X1TS U1280 ( .A(n2629), .B(\add_x_19_5/n42 ), .Y(n1408) );
  XNOR2X1TS U1281 ( .A(n1408), .B(\add_x_19_5/n43 ), .Y(
        \addr_calc/iir_write_addr[29] ) );
  OAI21X1TS U1282 ( .A0(\add_x_19_4/n154 ), .A1(\add_x_19_4/n156 ), .B0(
        \add_x_19_4/n155 ), .Y(n1409) );
  CLKINVX1TS U1283 ( .A(\add_x_19_4/n152 ), .Y(n1410) );
  OAI21XLTS U1284 ( .A0(\add_x_19_4/n151 ), .A1(n1410), .B0(n1409), .Y(n1411)
         );
  OAI31XLTS U1285 ( .A0(\add_x_19_4/n151 ), .A1(n1409), .A2(n1410), .B0(n1411), 
        .Y(\addr_calc/iir_read_addr[9] ) );
  OAI21X1TS U1286 ( .A0(\add_x_19_3/n165 ), .A1(\add_x_19_3/n167 ), .B0(
        \add_x_19_3/n166 ), .Y(n1412) );
  CLKINVX1TS U1287 ( .A(\add_x_19_3/n163 ), .Y(n1413) );
  OAI21XLTS U1288 ( .A0(\add_x_19_3/n162 ), .A1(n1413), .B0(n1412), .Y(n1414)
         );
  OAI31XLTS U1289 ( .A0(\add_x_19_3/n162 ), .A1(n1412), .A2(n1413), .B0(n1414), 
        .Y(\addr_calc/fir_write_addr[7] ) );
  NAND2X1TS U1290 ( .A(n2631), .B(\add_x_19_3/n42 ), .Y(n1415) );
  XNOR2X1TS U1291 ( .A(n1415), .B(\add_x_19_3/n43 ), .Y(
        \addr_calc/fir_write_addr[29] ) );
  NAND2X1TS U1292 ( .A(\add_x_19_2/n207 ), .B(\add_x_19_2/n111 ), .Y(n1416) );
  XNOR2X1TS U1293 ( .A(n1416), .B(\add_x_19_2/n112 ), .Y(
        \addr_calc/fir_read_addr[16] ) );
  OAI21XLTS U1294 ( .A0(\add_x_19_0/n154 ), .A1(\add_x_19_0/n156 ), .B0(
        \add_x_19_0/n155 ), .Y(n1417) );
  CLKINVX1TS U1295 ( .A(\add_x_19_0/n152 ), .Y(n1418) );
  OAI21XLTS U1296 ( .A0(\add_x_19_0/n151 ), .A1(n1418), .B0(n1417), .Y(n1419)
         );
  OAI31XLTS U1297 ( .A0(\add_x_19_0/n151 ), .A1(n1417), .A2(n1418), .B0(n1419), 
        .Y(\addr_calc/fft_read_addr[9] ) );
  NAND2X1TS U1298 ( .A(\add_x_19_0/n207 ), .B(\add_x_19_0/n111 ), .Y(n1420) );
  XNOR2X1TS U1299 ( .A(n1420), .B(\add_x_19_0/n112 ), .Y(
        \addr_calc/fft_read_addr[16] ) );
  NAND2BX1TS U1300 ( .AN(\add_x_19_2/n184 ), .B(\add_x_19_2/n185 ), .Y(n1421)
         );
  XOR2X1TS U1301 ( .A(\add_x_19_2/n186 ), .B(n1421), .Y(
        \addr_calc/fir_read_addr[2] ) );
  NAND2BX1TS U1302 ( .AN(\add_x_19_0/n188 ), .B(\add_x_19_0/n189 ), .Y(n1422)
         );
  XOR2X1TS U1303 ( .A(\add_x_19_0/n191 ), .B(n1422), .Y(
        \addr_calc/fft_read_addr[1] ) );
  CLKINVX1TS U1304 ( .A(\add_x_19_0/n182 ), .Y(n1423) );
  OAI21X1TS U1305 ( .A0(\add_x_19_0/n184 ), .A1(\add_x_19_0/n186 ), .B0(
        \add_x_19_0/n185 ), .Y(n1424) );
  OAI21XLTS U1306 ( .A0(\add_x_19_0/n181 ), .A1(n1423), .B0(n1424), .Y(n1425)
         );
  OAI31XLTS U1307 ( .A0(\add_x_19_0/n181 ), .A1(n1424), .A2(n1423), .B0(n1425), 
        .Y(\addr_calc/fft_read_addr[3] ) );
  OA21XLTS U1308 ( .A0(n2035), .A1(n2393), .B0(\add_x_19_1/n191 ), .Y(
        \addr_calc/fft_write_addr[0] ) );
  NAND4BX1TS U1309 ( .AN(\add_x_22_5/n35 ), .B(
        \addr_calc/iir_write_calc/count[23] ), .C(n2579), .D(\add_x_22_5/n43 ), 
        .Y(\add_x_22_5/n26 ) );
  NAND2BX1TS U1310 ( .AN(\add_x_22_0/n26 ), .B(\add_x_22_0/n59 ), .Y(
        \add_x_22_0/n24 ) );
  NAND3BX1TS U1311 ( .AN(\DP_OP_158_296_6262/n1792 ), .B(n1783), .C(
        \DP_OP_158_296_6262/n1837 ), .Y(\DP_OP_158_296_6262/n1834 ) );
  OAI21X1TS U1312 ( .A0(\add_x_19_5/n55 ), .A1(\add_x_19_5/n59 ), .B0(
        \add_x_19_5/n56 ), .Y(n1426) );
  AOI21X1TS U1313 ( .A0(\add_x_19_5/n53 ), .A1(\add_x_19_5/n62 ), .B0(n1426), 
        .Y(\add_x_19_5/n52 ) );
  NAND2BX1TS U1314 ( .AN(\add_x_22_5/n87 ), .B(\add_x_22_5/n93 ), .Y(
        \add_x_22_5/n85 ) );
  NAND2BX1TS U1315 ( .AN(\add_x_22_1/n87 ), .B(\add_x_22_1/n93 ), .Y(
        \add_x_22_1/n85 ) );
  NAND4BX1TS U1316 ( .AN(\add_x_22_3/n26 ), .B(\add_x_22_3/n59 ), .C(n1896), 
        .D(\add_x_22_3/n9 ), .Y(n1427) );
  NOR2BX1TS U1317 ( .AN(n1833), .B(n1427), .Y(\add_x_22_3/n2 ) );
  XNOR2X1TS U1318 ( .A(n1833), .B(n1427), .Y(
        \addr_calc/fir_write_calc/counter/N72 ) );
  NAND4BX1TS U1319 ( .AN(\add_x_22_4/n26 ), .B(\add_x_22_4/n59 ), .C(n2561), 
        .D(\add_x_22_4/n9 ), .Y(n1428) );
  NOR2BX1TS U1320 ( .AN(\addr_calc/iir_read_calc/count[29] ), .B(n1428), .Y(
        \add_x_22_4/n2 ) );
  XNOR2X1TS U1321 ( .A(\addr_calc/iir_read_calc/count[29] ), .B(n1428), .Y(
        \addr_calc/iir_read_calc/counter/N72 ) );
  NAND4BX1TS U1322 ( .AN(\add_x_22_2/n26 ), .B(\add_x_22_2/n59 ), .C(
        \addr_calc/fir_read_calc/count[28] ), .D(\add_x_22_2/n9 ), .Y(n1429)
         );
  NOR2BX1TS U1323 ( .AN(\addr_calc/fir_read_calc/count[29] ), .B(n1429), .Y(
        \add_x_22_2/n2 ) );
  XNOR2X1TS U1324 ( .A(\addr_calc/fir_read_calc/count[29] ), .B(n1429), .Y(
        \addr_calc/fir_read_calc/counter/N72 ) );
  NAND2BX1TS U1325 ( .AN(\add_x_19_1/n36 ), .B(\add_x_19_1/n37 ), .Y(n1430) );
  XOR2X1TS U1326 ( .A(\add_x_19_1/n38 ), .B(n1430), .Y(
        \addr_calc/fft_write_addr[30] ) );
  NAND2BX1TS U1327 ( .AN(\add_x_19_3/n100 ), .B(\add_x_19_3/n101 ), .Y(n1431)
         );
  XOR2X1TS U1328 ( .A(\add_x_19_3/n102 ), .B(n1431), .Y(
        \addr_calc/fir_write_addr[18] ) );
  NAND2BX1TS U1329 ( .AN(\add_x_19_2/n100 ), .B(\add_x_19_2/n101 ), .Y(n1432)
         );
  XOR2X1TS U1330 ( .A(\add_x_19_2/n102 ), .B(n1432), .Y(
        \addr_calc/fir_read_addr[18] ) );
  NAND2BX1TS U1331 ( .AN(\add_x_19_4/n81 ), .B(\add_x_19_4/n82 ), .Y(n1433) );
  NAND2BX1TS U1332 ( .AN(\add_x_19_0/n81 ), .B(\add_x_19_0/n82 ), .Y(n1434) );
  XOR2X1TS U1333 ( .A(\add_x_19_0/n83 ), .B(n1434), .Y(
        \addr_calc/fft_read_addr[22] ) );
  NAND2BX1TS U1334 ( .AN(\add_x_19_3/n58 ), .B(\add_x_19_3/n59 ), .Y(n1435) );
  XOR2X1TS U1335 ( .A(\add_x_19_3/n60 ), .B(n1435), .Y(
        \addr_calc/fir_write_addr[26] ) );
  NAND2BX1TS U1336 ( .AN(\add_x_19_5/n165 ), .B(\add_x_19_5/n166 ), .Y(n1436)
         );
  XOR2X1TS U1337 ( .A(\add_x_19_5/n167 ), .B(n1436), .Y(
        \addr_calc/iir_write_addr[6] ) );
  NAND2BX1TS U1338 ( .AN(\add_x_19_4/n131 ), .B(\add_x_19_4/n132 ), .Y(n1437)
         );
  XOR2X1TS U1339 ( .A(\add_x_19_4/n133 ), .B(n1437), .Y(
        \addr_calc/iir_read_addr[12] ) );
  NAND2BX1TS U1340 ( .AN(\add_x_19_3/n89 ), .B(\add_x_19_3/n90 ), .Y(n1438) );
  XOR2X1TS U1341 ( .A(\add_x_19_3/n91 ), .B(n1438), .Y(
        \addr_calc/fir_write_addr[20] ) );
  NAND2BX1TS U1342 ( .AN(\add_x_19_2/n123 ), .B(\add_x_19_2/n124 ), .Y(n1439)
         );
  XOR2X1TS U1343 ( .A(\add_x_19_2/n125 ), .B(n1439), .Y(
        \addr_calc/fir_read_addr[14] ) );
  NAND2BX1TS U1344 ( .AN(\add_x_19_1/n131 ), .B(\add_x_19_1/n132 ), .Y(n1440)
         );
  XOR2X1TS U1345 ( .A(\add_x_19_1/n133 ), .B(n1440), .Y(
        \addr_calc/fft_write_addr[12] ) );
  NAND2BX1TS U1346 ( .AN(\add_x_19_1/n89 ), .B(\add_x_19_1/n90 ), .Y(n1441) );
  NAND2BX1TS U1347 ( .AN(\add_x_19_0/n123 ), .B(\add_x_19_0/n124 ), .Y(n1442)
         );
  XOR2X1TS U1348 ( .A(\add_x_19_0/n125 ), .B(n1442), .Y(
        \addr_calc/fft_read_addr[14] ) );
  NAND2X1TS U1349 ( .A(\add_x_19_4/n207 ), .B(\add_x_19_4/n111 ), .Y(n1443) );
  XNOR2X1TS U1350 ( .A(n1443), .B(\add_x_19_4/n112 ), .Y(
        \addr_calc/iir_read_addr[16] ) );
  NAND2X1TS U1351 ( .A(\add_x_19_2/n213 ), .B(\add_x_19_2/n145 ), .Y(n1444) );
  XNOR2X1TS U1352 ( .A(n1444), .B(\add_x_19_2/n146 ), .Y(
        \addr_calc/fir_read_addr[10] ) );
  NAND2X1TS U1353 ( .A(n2633), .B(\add_x_19_2/n42 ), .Y(n1445) );
  XNOR2X1TS U1354 ( .A(n1445), .B(\add_x_19_2/n43 ), .Y(
        \addr_calc/fir_read_addr[29] ) );
  NAND2X1TS U1355 ( .A(\add_x_19_1/n213 ), .B(\add_x_19_1/n145 ), .Y(n1446) );
  NAND2X1TS U1356 ( .A(\add_x_19_1/n207 ), .B(\add_x_19_1/n111 ), .Y(n1447) );
  OAI21X1TS U1357 ( .A0(\add_x_19_0/n165 ), .A1(\add_x_19_0/n167 ), .B0(
        \add_x_19_0/n166 ), .Y(n1448) );
  CLKINVX1TS U1358 ( .A(\add_x_19_0/n163 ), .Y(n1449) );
  OAI21X1TS U1359 ( .A0(\add_x_19_0/n162 ), .A1(n1449), .B0(n1448), .Y(n1450)
         );
  OAI31X1TS U1360 ( .A0(\add_x_19_0/n162 ), .A1(n1448), .A2(n1449), .B0(n1450), 
        .Y(\addr_calc/fft_read_addr[7] ) );
  NAND2X1TS U1361 ( .A(n2628), .B(\add_x_19_0/n42 ), .Y(n1451) );
  XNOR2X1TS U1362 ( .A(n1451), .B(\add_x_19_0/n43 ), .Y(
        \addr_calc/fft_read_addr[29] ) );
  NAND3X1TS U1363 ( .A(n802), .B(n2310), .C(n2055), .Y(n1452) );
  AOI211X1TS U1364 ( .A0(n2336), .A1(n2311), .B0(acc_done), .C0(n1452), .Y(
        \pla_top/N59 ) );
  NAND2BX1TS U1365 ( .AN(\add_x_19_1/n188 ), .B(\add_x_19_1/n189 ), .Y(n1453)
         );
  XOR2X1TS U1366 ( .A(\add_x_19_1/n191 ), .B(n1453), .Y(
        \addr_calc/fft_write_addr[1] ) );
  NAND2BX1TS U1367 ( .AN(\add_x_19_1/n184 ), .B(\add_x_19_1/n185 ), .Y(n1454)
         );
  XOR2X1TS U1368 ( .A(\add_x_19_1/n186 ), .B(n1454), .Y(
        \addr_calc/fft_write_addr[2] ) );
  OA21XLTS U1369 ( .A0(\addr_calc/fft_read_calc/count[0] ), .A1(n2393), .B0(
        \add_x_19_0/n191 ), .Y(\addr_calc/fft_read_addr[0] ) );
  NOR3BX1TS U1370 ( .AN(n936), .B(data_to_fir), .C(\data_cntl/N95 ), .Y(
        \data_cntl/N264 ) );
  XOR2X4TS U1371 ( .A(n1661), .B(\add_x_22_4/n15 ), .Y(
        \DP_OP_159_297_3515/n87 ) );
  XOR2X4TS U1372 ( .A(\DP_OP_158_296_6262/n1998 ), .B(n2366), .Y(n2593) );
  XOR2X4TS U1373 ( .A(\DP_OP_159_297_3515/n792 ), .B(n1964), .Y(
        \DP_OP_159_297_3515/n556 ) );
  XNOR2X4TS U1374 ( .A(n1568), .B(n1569), .Y(\addr_calc/fir_read_addr[21] ) );
  NOR2XLTS U1375 ( .A(\DP_OP_158_296_6262/n1891 ), .B(n1515), .Y(
        \DP_OP_158_296_6262/n1883 ) );
  NAND2X2TS U1376 ( .A(\DP_OP_159_297_3515/n648 ), .B(
        \DP_OP_159_297_3515/n672 ), .Y(\DP_OP_159_297_3515/n646 ) );
  XNOR2X4TS U1377 ( .A(n2617), .B(n2570), .Y(\DP_OP_159_297_3515/n674 ) );
  NOR2X4TS U1378 ( .A(\DP_OP_159_297_3515/n102 ), .B(\DP_OP_159_297_3515/n87 ), 
        .Y(\DP_OP_159_297_3515/n85 ) );
  XOR2X4TS U1379 ( .A(n1738), .B(n2033), .Y(\DP_OP_159_297_3515/n116 ) );
  NAND2XLTS U1380 ( .A(\addr_calc/iir_read_calc/count[2] ), .B(n2444), .Y(
        \add_x_19_4/n185 ) );
  AO22X2TS U1381 ( .A0(n1714), .A1(\addr_calc/iir_read_calc/counter/N50 ), 
        .B0(n2648), .B1(n1905), .Y(n964) );
  XNOR2X2TS U1382 ( .A(\add_x_19_1/n65 ), .B(\add_x_19_1/n7 ), .Y(
        \addr_calc/fft_write_addr[25] ) );
  XNOR2X2TS U1383 ( .A(\add_x_19_1/n50 ), .B(\add_x_19_1/n4 ), .Y(
        \addr_calc/fft_write_addr[28] ) );
  NOR2X2TS U1384 ( .A(\DP_OP_158_296_6262/n277 ), .B(\DP_OP_158_296_6262/n266 ), .Y(\DP_OP_158_296_6262/n264 ) );
  XOR2X4TS U1385 ( .A(n1655), .B(n1946), .Y(\DP_OP_158_296_6262/n998 ) );
  NAND2X2TS U1386 ( .A(\DP_OP_159_297_3515/n1024 ), .B(
        \DP_OP_159_297_3515/n873 ), .Y(n1734) );
  NAND2X4TS U1387 ( .A(n1788), .B(\DP_OP_159_297_3515/n1025 ), .Y(
        \DP_OP_159_297_3515/n1024 ) );
  INVX4TS U1388 ( .A(n1786), .Y(n1787) );
  INVXLTS U1389 ( .A(\DP_OP_158_296_6262/n1959 ), .Y(n1455) );
  XNOR2X2TS U1390 ( .A(\add_x_19_2/n122 ), .B(\add_x_19_2/n17 ), .Y(
        \addr_calc/fir_read_addr[15] ) );
  XOR2X2TS U1391 ( .A(\DP_OP_159_297_3515/n1057 ), .B(
        \DP_OP_159_297_3515/n878 ), .Y(n2610) );
  NOR2X2TS U1392 ( .A(\DP_OP_159_297_3515/n1063 ), .B(
        \DP_OP_159_297_3515/n879 ), .Y(\DP_OP_159_297_3515/n1057 ) );
  OAI21X2TS U1393 ( .A0(\add_x_19_2/n83 ), .A1(\add_x_19_2/n81 ), .B0(
        \add_x_19_2/n82 ), .Y(n1596) );
  INVX6TS U1394 ( .A(n1786), .Y(n1788) );
  CLKBUFX2TS U1395 ( .A(n1641), .Y(n1456) );
  NAND2X4TS U1396 ( .A(n1624), .B(n1623), .Y(\DP_OP_159_297_3515/n18 ) );
  XNOR2X2TS U1397 ( .A(n1756), .B(n2046), .Y(\DP_OP_158_296_6262/n1171 ) );
  NAND2X2TS U1398 ( .A(n1511), .B(n1501), .Y(\DP_OP_159_297_3515/n1026 ) );
  AOI21X4TS U1399 ( .A0(\add_x_19_1/n43 ), .A1(n2632), .B0(n1546), .Y(
        \add_x_19_1/n38 ) );
  INVX2TS U1400 ( .A(n2419), .Y(n2421) );
  NOR2X4TS U1401 ( .A(n1501), .B(n1487), .Y(n1591) );
  INVX2TS U1402 ( .A(n1486), .Y(n1487) );
  AO22X4TS U1403 ( .A0(n1769), .A1(\addr_calc/iir_write_calc/counter/N64 ), 
        .B0(n2672), .B1(\addr_calc/iir_write_calc/count[21] ), .Y(n981) );
  XNOR2X1TS U1404 ( .A(n2608), .B(n2562), .Y(\DP_OP_159_297_3515/n723 ) );
  XOR2X4TS U1405 ( .A(n1787), .B(\DP_OP_159_297_3515/n875 ), .Y(n2608) );
  NAND2X2TS U1406 ( .A(n1831), .B(n1503), .Y(\DP_OP_159_297_3515/n998 ) );
  INVX2TS U1407 ( .A(n1502), .Y(n1503) );
  XOR2X2TS U1408 ( .A(\DP_OP_158_296_6262/n829 ), .B(n1838), .Y(n1653) );
  NOR2X4TS U1409 ( .A(n1693), .B(\DP_OP_158_296_6262/n1951 ), .Y(
        \DP_OP_158_296_6262/n1950 ) );
  INVX2TS U1410 ( .A(n1513), .Y(\DP_OP_158_296_6262/n1952 ) );
  INVX2TS U1411 ( .A(n1501), .Y(\DP_OP_158_296_6262/n1966 ) );
  INVX2TS U1412 ( .A(n1500), .Y(n1501) );
  NOR2X4TS U1413 ( .A(n1485), .B(n1815), .Y(\DP_OP_158_296_6262/n1862 ) );
  NOR2X4TS U1414 ( .A(n1794), .B(\DP_OP_158_296_6262/n1841 ), .Y(
        \DP_OP_158_296_6262/n1840 ) );
  XNOR2X4TS U1415 ( .A(n1463), .B(\addr_calc/fft_read_calc/count[29] ), .Y(
        \DP_OP_158_296_6262/n933 ) );
  INVX2TS U1416 ( .A(n1483), .Y(n1485) );
  CLKINVX3TS U1417 ( .A(filesize[2]), .Y(n1641) );
  OAI21X2TS U1418 ( .A0(\add_x_19_2/n44 ), .A1(\add_x_19_2/n113 ), .B0(
        \add_x_19_2/n45 ), .Y(\add_x_19_2/n43 ) );
  INVX2TS U1419 ( .A(n1481), .Y(n1482) );
  INVX4TS U1420 ( .A(\DP_OP_158_296_6262/n2048 ), .Y(\DP_OP_158_296_6262/n841 ) );
  XNOR2X2TS U1421 ( .A(\DP_OP_158_296_6262/n2048 ), .B(\add_x_22_0/n49 ), .Y(
        n1459) );
  CLKINVX3TS U1422 ( .A(n2787), .Y(n1458) );
  INVX2TS U1423 ( .A(n1746), .Y(n1673) );
  NOR2X4TS U1424 ( .A(n1459), .B(\DP_OP_158_296_6262/n1079 ), .Y(
        \DP_OP_158_296_6262/n1077 ) );
  AO22X4TS U1425 ( .A0(n1152), .A1(\addr_calc/fir_write_calc/counter/N52 ), 
        .B0(n1261), .B1(n1872), .Y(n1121) );
  BUFX8TS U1426 ( .A(n2671), .Y(n2662) );
  OAI2BB1X2TS U1427 ( .A0N(n2009), .A1N(n1263), .B0(n1618), .Y(n1110) );
  XOR2X4TS U1428 ( .A(\DP_OP_159_297_3515/n892 ), .B(n2341), .Y(n2625) );
  CLKINVX6TS U1429 ( .A(\addr_calc/fft_read_calc/counter/N38 ), .Y(n783) );
  XOR2X4TS U1430 ( .A(n1149), .B(n1943), .Y(\DP_OP_158_296_6262/n962 ) );
  NOR2X6TS U1431 ( .A(n1696), .B(n1461), .Y(n2807) );
  XNOR2X2TS U1432 ( .A(n1149), .B(n1873), .Y(\DP_OP_158_296_6262/n68 ) );
  INVX4TS U1433 ( .A(n1742), .Y(n1743) );
  INVX2TS U1434 ( .A(n1742), .Y(n1672) );
  INVX2TS U1435 ( .A(n1742), .Y(n1744) );
  CLKINVX6TS U1436 ( .A(n1741), .Y(n1745) );
  AND2X8TS U1437 ( .A(n1716), .B(n1715), .Y(n1461) );
  NOR2X4TS U1438 ( .A(n1796), .B(\DP_OP_158_296_6262/n1882 ), .Y(
        \DP_OP_158_296_6262/n1881 ) );
  XOR2X4TS U1439 ( .A(\DP_OP_159_297_3515/n792 ), .B(\add_x_22_4/n30 ), .Y(
        \DP_OP_159_297_3515/n131 ) );
  AO22X2TS U1440 ( .A0(n1151), .A1(\addr_calc/fir_read_calc/counter/N53 ), 
        .B0(\addr_calc/fir_read_calc/count[10] ), .B1(n1741), .Y(n1088) );
  AO22X2TS U1441 ( .A0(n1821), .A1(\addr_calc/fir_read_calc/counter/N64 ), 
        .B0(\addr_calc/fir_read_calc/count[21] ), .B1(n1741), .Y(n1077) );
  NOR2X4TS U1442 ( .A(\DP_OP_158_296_6262/n1111 ), .B(
        \DP_OP_158_296_6262/n1124 ), .Y(\DP_OP_158_296_6262/n1109 ) );
  XNOR2X4TS U1443 ( .A(n1729), .B(n1960), .Y(\DP_OP_158_296_6262/n1111 ) );
  NAND2X2TS U1444 ( .A(\add_x_22_1/n4 ), .B(\add_x_22_1/n59 ), .Y(
        \add_x_22_1/n3 ) );
  XNOR2X1TS U1445 ( .A(n1871), .B(n1775), .Y(\DP_OP_158_296_6262/n54 ) );
  OAI21X2TS U1446 ( .A0(\add_x_19_2/n156 ), .A1(\add_x_19_2/n135 ), .B0(
        \add_x_19_2/n136 ), .Y(\add_x_19_2/n134 ) );
  NOR2X4TS U1447 ( .A(n1693), .B(\DP_OP_158_296_6262/n1965 ), .Y(
        \DP_OP_158_296_6262/n1964 ) );
  AND2X8TS U1448 ( .A(\DP_OP_158_296_6262/n1791 ), .B(
        \DP_OP_158_296_6262/n1869 ), .Y(n1462) );
  INVX6TS U1449 ( .A(n1677), .Y(n1717) );
  AO22X4TS U1450 ( .A0(n1712), .A1(\addr_calc/iir_read_calc/counter/N60 ), 
        .B0(n2650), .B1(\addr_calc/iir_read_calc/count[17] ), .Y(n954) );
  XNOR2X2TS U1451 ( .A(\add_x_19_1/n122 ), .B(\add_x_19_1/n17 ), .Y(
        \addr_calc/fft_write_addr[15] ) );
  XNOR2X2TS U1452 ( .A(n1652), .B(\addr_calc/fir_read_calc/count[22] ), .Y(
        \DP_OP_158_296_6262/n148 ) );
  AO22X4TS U1453 ( .A0(n1721), .A1(\addr_calc/fft_write_calc/counter/N60 ), 
        .B0(n2667), .B1(n1924), .Y(n1049) );
  AO22X4TS U1454 ( .A0(n1724), .A1(\addr_calc/fft_write_calc/counter/N59 ), 
        .B0(n2666), .B1(n2567), .Y(n1050) );
  XOR2X2TS U1455 ( .A(\DP_OP_158_296_6262/n829 ), .B(n1859), .Y(n1471) );
  NOR2X8TS U1456 ( .A(n1795), .B(\DP_OP_158_296_6262/n1848 ), .Y(
        \DP_OP_158_296_6262/n1847 ) );
  XOR2X4TS U1457 ( .A(\DP_OP_158_296_6262/n1840 ), .B(n1464), .Y(n1463) );
  NOR2X4TS U1458 ( .A(\DP_OP_158_296_6262/n1903 ), .B(
        \DP_OP_158_296_6262/n1877 ), .Y(\DP_OP_158_296_6262/n1791 ) );
  NAND2X4TS U1459 ( .A(\DP_OP_158_296_6262/n1890 ), .B(
        \DP_OP_158_296_6262/n1878 ), .Y(\DP_OP_158_296_6262/n1877 ) );
  NAND2X2TS U1460 ( .A(\DP_OP_158_296_6262/n1791 ), .B(
        \DP_OP_158_296_6262/n1849 ), .Y(\DP_OP_158_296_6262/n1848 ) );
  AO22X4TS U1461 ( .A0(n1727), .A1(\addr_calc/fft_write_calc/counter/N48 ), 
        .B0(n2663), .B1(n1479), .Y(n1061) );
  XOR2X4TS U1462 ( .A(\DP_OP_158_296_6262/n1840 ), .B(n1464), .Y(n1777) );
  XNOR2X4TS U1463 ( .A(\add_x_19_1/n80 ), .B(\add_x_19_1/n9 ), .Y(
        \addr_calc/fft_write_addr[23] ) );
  OR2X4TS U1464 ( .A(\DP_OP_158_296_6262/n2011 ), .B(
        \DP_OP_158_296_6262/n1987 ), .Y(n1693) );
  INVX2TS U1465 ( .A(n1506), .Y(\DP_OP_159_297_3515/n876 ) );
  XNOR2X4TS U1466 ( .A(n2615), .B(n1951), .Y(\DP_OP_159_297_3515/n650 ) );
  NOR2X4TS U1467 ( .A(\addr_calc/fir_read_calc/count[7] ), .B(n2421), .Y(
        \add_x_19_2/n162 ) );
  NAND2X2TS U1468 ( .A(\addr_calc/fir_read_calc/count[7] ), .B(n2421), .Y(
        \add_x_19_2/n163 ) );
  XNOR2X4TS U1469 ( .A(\add_x_19_2/n35 ), .B(\add_x_19_2/n1 ), .Y(
        \addr_calc/fir_read_addr[31] ) );
  INVX2TS U1470 ( .A(n1514), .Y(n1516) );
  NAND2X4TS U1471 ( .A(\DP_OP_158_296_6262/n960 ), .B(
        \DP_OP_158_296_6262/n996 ), .Y(\DP_OP_158_296_6262/n958 ) );
  NOR2X2TS U1472 ( .A(\DP_OP_158_296_6262/n1896 ), .B(n2589), .Y(
        \DP_OP_158_296_6262/n1895 ) );
  NOR2X4TS U1473 ( .A(\DP_OP_158_296_6262/n129 ), .B(\DP_OP_158_296_6262/n64 ), 
        .Y(\DP_OP_158_296_6262/n62 ) );
  NOR2X4TS U1474 ( .A(n1717), .B(\DP_OP_158_296_6262/n1854 ), .Y(n1736) );
  INVX8TS U1475 ( .A(n1793), .Y(n1795) );
  AOI21X2TS U1476 ( .A0(\add_x_19_2/n69 ), .A1(\add_x_19_2/n61 ), .B0(
        \add_x_19_2/n62 ), .Y(\add_x_19_2/n60 ) );
  OAI21X2TS U1477 ( .A0(\add_x_19_2/n113 ), .A1(\add_x_19_2/n93 ), .B0(
        \add_x_19_2/n94 ), .Y(\add_x_19_2/n92 ) );
  NOR2X4TS U1478 ( .A(\DP_OP_158_296_6262/n1023 ), .B(
        \DP_OP_158_296_6262/n958 ), .Y(\DP_OP_158_296_6262/n956 ) );
  NAND2X4TS U1479 ( .A(\DP_OP_158_296_6262/n1025 ), .B(
        \DP_OP_158_296_6262/n1053 ), .Y(\DP_OP_158_296_6262/n1023 ) );
  INVX6TS U1480 ( .A(n1793), .Y(n1794) );
  NOR2X4TS U1481 ( .A(n1794), .B(\DP_OP_158_296_6262/n1861 ), .Y(
        \DP_OP_158_296_6262/n1860 ) );
  INVX2TS U1482 ( .A(n1492), .Y(n1493) );
  OAI2BB2X2TS U1483 ( .B0(n1740), .B1(\add_x_22_5/n71 ), .A0N(n1773), .A1N(
        \addr_calc/iir_write_calc/counter/N56 ), .Y(n989) );
  XNOR2X4TS U1484 ( .A(n2621), .B(n1940), .Y(\DP_OP_159_297_3515/n714 ) );
  INVX2TS U1485 ( .A(n1496), .Y(n1497) );
  INVX6TS U1486 ( .A(n2661), .Y(n1474) );
  XOR2X4TS U1487 ( .A(n1796), .B(n2361), .Y(n2594) );
  INVX2TS U1488 ( .A(n1519), .Y(n1520) );
  XNOR2X4TS U1489 ( .A(\add_x_19_1/n57 ), .B(\add_x_19_1/n5 ), .Y(
        \addr_calc/fft_write_addr[27] ) );
  NOR2X4TS U1490 ( .A(n1499), .B(n1491), .Y(\DP_OP_158_296_6262/n1890 ) );
  INVX2TS U1491 ( .A(n1490), .Y(n1491) );
  INVX2TS U1492 ( .A(n1498), .Y(n1499) );
  NOR2X4TS U1493 ( .A(n1795), .B(\DP_OP_158_296_6262/n1903 ), .Y(n1642) );
  INVX2TS U1494 ( .A(n1488), .Y(n1489) );
  NOR2X2TS U1495 ( .A(n1505), .B(n1510), .Y(\DP_OP_158_296_6262/n1973 ) );
  INVXLTS U1496 ( .A(\DP_OP_158_296_6262/n1945 ), .Y(
        \DP_OP_158_296_6262/n1946 ) );
  BUFX8TS U1497 ( .A(n2797), .Y(n2671) );
  INVX2TS U1498 ( .A(n2005), .Y(n2006) );
  INVX2TS U1499 ( .A(n1523), .Y(\DP_OP_158_296_6262/n1911 ) );
  INVX2TS U1500 ( .A(n1814), .Y(n1815) );
  CLKINVX3TS U1501 ( .A(n1917), .Y(n1918) );
  INVX2TS U1502 ( .A(\addr_calc/fir_write_calc/count[2] ), .Y(n1989) );
  INVX2TS U1503 ( .A(\addr_calc/fft_read_calc/count[0] ), .Y(n2057) );
  INVX2TS U1504 ( .A(n1807), .Y(n2330) );
  INVX2TS U1505 ( .A(\add_x_19_5/n36 ), .Y(n1533) );
  AND2X2TS U1506 ( .A(\add_x_19_0/n196 ), .B(\add_x_19_0/n56 ), .Y(n1465) );
  AND2X2TS U1507 ( .A(\add_x_19_4/n200 ), .B(\add_x_19_4/n79 ), .Y(n1466) );
  INVXLTS U1508 ( .A(n1521), .Y(\DP_OP_159_297_3515/n869 ) );
  AND2X2TS U1509 ( .A(\add_x_19_4/n199 ), .B(\add_x_19_4/n67 ), .Y(n1467) );
  OR3X1TS U1510 ( .A(\data_cntl/N159 ), .B(n2790), .C(n1861), .Y(n1468) );
  INVX4TS U1511 ( .A(n1959), .Y(n1960) );
  INVX2TS U1512 ( .A(n1815), .Y(\DP_OP_158_296_6262/n1869 ) );
  INVXLTS U1513 ( .A(\DP_OP_158_296_6262/n1966 ), .Y(n2367) );
  INVXLTS U1514 ( .A(n1831), .Y(\DP_OP_159_297_3515/n870 ) );
  INVXLTS U1515 ( .A(\DP_OP_158_296_6262/n1952 ), .Y(n2368) );
  INVX4TS U1516 ( .A(n1677), .Y(n1796) );
  CLKINVX6TS U1517 ( .A(n2589), .Y(n1677) );
  XNOR2X4TS U1518 ( .A(\DP_OP_158_296_6262/n1978 ), .B(n2365), .Y(n1469) );
  INVX2TS U1519 ( .A(n1545), .Y(\add_x_19_3/n123 ) );
  AND2X2TS U1520 ( .A(\add_x_19_3/n72 ), .B(\add_x_19_3/n46 ), .Y(n1470) );
  INVXLTS U1521 ( .A(\DP_OP_159_297_3515/n880 ), .Y(n2371) );
  INVXLTS U1522 ( .A(n1817), .Y(n2370) );
  BUFX6TS U1523 ( .A(n2680), .Y(n2673) );
  INVX2TS U1524 ( .A(\addr_calc/iir_read_calc/count[3] ), .Y(n1901) );
  INVX2TS U1525 ( .A(\addr_calc/iir_read_calc/count[25] ), .Y(n1925) );
  INVX2TS U1526 ( .A(\addr_calc/fft_write_calc/count[6] ), .Y(n2029) );
  INVX2TS U1527 ( .A(\addr_calc/fir_read_calc/count[10] ), .Y(n1897) );
  INVX2TS U1528 ( .A(n1986), .Y(\addr_calc/fir_write_calc/counter/N43 ) );
  CLKBUFX2TS U1529 ( .A(\add_x_19_5/n59 ), .Y(n1473) );
  CLKINVX3TS U1530 ( .A(n1474), .Y(n1476) );
  CLKBUFX2TS U1531 ( .A(\addr_calc/fir_read_calc/count[7] ), .Y(n1480) );
  INVXLTS U1532 ( .A(filesize[14]), .Y(n1481) );
  INVXLTS U1533 ( .A(filesize[25]), .Y(n1483) );
  INVXLTS U1534 ( .A(n1483), .Y(n1484) );
  INVXLTS U1535 ( .A(filesize[11]), .Y(n1486) );
  INVXLTS U1536 ( .A(filesize[7]), .Y(n1488) );
  INVXLTS U1537 ( .A(filesize[20]), .Y(n1490) );
  INVXLTS U1538 ( .A(filesize[5]), .Y(n1492) );
  INVXLTS U1539 ( .A(filesize[6]), .Y(n1494) );
  INVXLTS U1540 ( .A(filesize[4]), .Y(n1496) );
  INVXLTS U1541 ( .A(filesize[21]), .Y(n1498) );
  INVXLTS U1542 ( .A(filesize[10]), .Y(n1500) );
  INVXLTS U1543 ( .A(filesize[13]), .Y(n1502) );
  INVXLTS U1544 ( .A(filesize[8]), .Y(n1504) );
  INVXLTS U1545 ( .A(filesize[26]), .Y(n1507) );
  INVX2TS U1546 ( .A(n1507), .Y(n1508) );
  INVXLTS U1547 ( .A(filesize[9]), .Y(n1509) );
  INVXLTS U1548 ( .A(filesize[12]), .Y(n1512) );
  INVXLTS U1549 ( .A(filesize[22]), .Y(n1514) );
  INVXLTS U1550 ( .A(n1514), .Y(n1515) );
  INVXLTS U1551 ( .A(filesize[23]), .Y(n1517) );
  INVXLTS U1552 ( .A(filesize[15]), .Y(n1519) );
  INVXLTS U1553 ( .A(n1519), .Y(n1521) );
  INVXLTS U1554 ( .A(filesize[18]), .Y(n1522) );
  INVX2TS U1555 ( .A(n1522), .Y(n1523) );
  INVXLTS U1556 ( .A(filesize[0]), .Y(n1524) );
  INVX2TS U1557 ( .A(n1524), .Y(n1525) );
  INVXLTS U1558 ( .A(filesize[3]), .Y(n1526) );
  INVXLTS U1559 ( .A(filesize[16]), .Y(n1528) );
  INVX2TS U1560 ( .A(n1528), .Y(n1529) );
  NAND2X1TS U1561 ( .A(n1495), .B(n1493), .Y(\DP_OP_159_297_3515/n1052 ) );
  INVXLTS U1562 ( .A(n1495), .Y(\DP_OP_159_297_3515/n878 ) );
  INVXLTS U1563 ( .A(n1499), .Y(\DP_OP_159_297_3515/n950 ) );
  NAND2X1TS U1564 ( .A(n1499), .B(n1515), .Y(\DP_OP_159_297_3515/n943 ) );
  INVXLTS U1565 ( .A(filesize[19]), .Y(n1530) );
  INVX2TS U1566 ( .A(n1530), .Y(n1531) );
  AOI21X1TS U1567 ( .A0(\add_x_19_4/n134 ), .A1(\add_x_19_4/n126 ), .B0(
        \add_x_19_4/n127 ), .Y(\add_x_19_4/n125 ) );
  OAI21X1TS U1568 ( .A0(\add_x_19_5/n125 ), .A1(\add_x_19_5/n123 ), .B0(
        \add_x_19_5/n124 ), .Y(n1536) );
  OAI21X2TS U1569 ( .A0(\add_x_19_2/n38 ), .A1(\add_x_19_2/n36 ), .B0(
        \add_x_19_2/n37 ), .Y(\add_x_19_2/n35 ) );
  CLKINVX1TS U1570 ( .A(\add_x_19_1/n78 ), .Y(\add_x_19_1/n200 ) );
  AO21X4TS U1571 ( .A0(n1532), .A1(\add_x_19_5/n43 ), .B0(n1534), .Y(
        \add_x_19_5/n35 ) );
  XNOR2X2TS U1572 ( .A(\add_x_19_5/n35 ), .B(\add_x_19_5/n1 ), .Y(
        \addr_calc/iir_write_addr[31] ) );
  OAI21X1TS U1573 ( .A0(\add_x_19_5/n94 ), .A1(\add_x_19_5/n74 ), .B0(
        \add_x_19_5/n75 ), .Y(\add_x_19_5/n73 ) );
  NAND2X2TS U1574 ( .A(n2046), .B(n2409), .Y(\add_x_19_0/n132 ) );
  AOI21X1TS U1575 ( .A0(\add_x_19_5/n73 ), .A1(\add_x_19_5/n46 ), .B0(
        \add_x_19_5/n47 ), .Y(\add_x_19_5/n45 ) );
  NAND2X1TS U1576 ( .A(\add_x_19_5/n72 ), .B(\add_x_19_5/n46 ), .Y(
        \add_x_19_5/n44 ) );
  OAI21X2TS U1577 ( .A0(\add_x_19_5/n113 ), .A1(\add_x_19_5/n44 ), .B0(
        \add_x_19_5/n45 ), .Y(\add_x_19_5/n43 ) );
  OAI21X2TS U1578 ( .A0(\add_x_19_5/n156 ), .A1(\add_x_19_5/n135 ), .B0(
        \add_x_19_5/n136 ), .Y(\add_x_19_5/n134 ) );
  AOI21X4TS U1579 ( .A0(\add_x_19_3/n43 ), .A1(n2631), .B0(n1535), .Y(
        \add_x_19_3/n38 ) );
  XNOR2X2TS U1580 ( .A(n1536), .B(n1537), .Y(\addr_calc/iir_write_addr[15] )
         );
  INVX1TS U1581 ( .A(n1480), .Y(\add_x_22_2/n98 ) );
  CLKINVX1TS U1582 ( .A(\add_x_19_2/n162 ), .Y(\add_x_19_2/n216 ) );
  INVX2TS U1583 ( .A(\add_x_19_2/n157 ), .Y(\add_x_19_2/n156 ) );
  OAI21X2TS U1584 ( .A0(n1539), .A1(\add_x_19_0/n136 ), .B0(\add_x_19_0/n117 ), 
        .Y(\add_x_19_0/n115 ) );
  NOR2X2TS U1585 ( .A(n1539), .B(\add_x_19_0/n135 ), .Y(\add_x_19_0/n114 ) );
  NAND2X2TS U1586 ( .A(\add_x_19_0/n118 ), .B(\add_x_19_0/n126 ), .Y(n1539) );
  NAND2X1TS U1587 ( .A(\addr_calc/fir_write_calc/count[0] ), .B(n2393), .Y(
        \add_x_19_3/n191 ) );
  NAND2X2TS U1588 ( .A(n1990), .B(n2444), .Y(\add_x_19_3/n185 ) );
  NOR2X2TS U1589 ( .A(n1540), .B(n2413), .Y(\add_x_19_2/n144 ) );
  NAND2X2TS U1590 ( .A(n1540), .B(n2414), .Y(\add_x_19_2/n145 ) );
  XNOR2XLTS U1591 ( .A(n1656), .B(n1540), .Y(\DP_OP_158_296_6262/n297 ) );
  INVX1TS U1592 ( .A(\add_x_19_2/n145 ), .Y(\add_x_19_2/n143 ) );
  INVX2TS U1593 ( .A(\add_x_19_2/n113 ), .Y(\add_x_19_2/n112 ) );
  AOI21X2TS U1594 ( .A0(\add_x_19_2/n43 ), .A1(n2633), .B0(n1559), .Y(
        \add_x_19_2/n38 ) );
  XNOR2X1TS U1595 ( .A(\add_x_22_0/n1 ), .B(n1856), .Y(n1543) );
  OAI2BB1X1TS U1596 ( .A0N(\addr_calc/fft_read_calc/count[31] ), .A1N(n2658), 
        .B0(n1542), .Y(n1035) );
  XNOR2X1TS U1597 ( .A(\add_x_19_0/n38 ), .B(n1544), .Y(
        \addr_calc/fft_read_addr[30] ) );
  OAI21X1TS U1598 ( .A0(\add_x_19_3/n176 ), .A1(\add_x_19_3/n170 ), .B0(
        \add_x_19_3/n171 ), .Y(\add_x_19_3/n169 ) );
  AOI21X2TS U1599 ( .A0(\add_x_19_4/n179 ), .A1(\add_x_19_4/n187 ), .B0(
        \add_x_19_4/n180 ), .Y(\add_x_19_4/n178 ) );
  OAI21X1TS U1600 ( .A0(\add_x_19_3/n191 ), .A1(\add_x_19_3/n188 ), .B0(
        \add_x_19_3/n189 ), .Y(\add_x_19_3/n187 ) );
  OAI21X2TS U1601 ( .A0(\add_x_19_2/n151 ), .A1(\add_x_19_2/n155 ), .B0(
        \add_x_19_2/n152 ), .Y(\add_x_19_2/n150 ) );
  AOI21X1TS U1602 ( .A0(\add_x_19_2/n73 ), .A1(\add_x_19_2/n46 ), .B0(
        \add_x_19_2/n47 ), .Y(\add_x_19_2/n45 ) );
  NAND2X1TS U1603 ( .A(\add_x_19_5/n118 ), .B(\add_x_19_5/n126 ), .Y(
        \add_x_19_5/n116 ) );
  NOR2X1TS U1604 ( .A(\add_x_19_2/n181 ), .B(\add_x_19_2/n184 ), .Y(n1547) );
  AOI21X2TS U1605 ( .A0(n1547), .A1(\add_x_19_2/n187 ), .B0(n1548), .Y(
        \add_x_19_2/n178 ) );
  OAI21X1TS U1606 ( .A0(\add_x_19_5/n136 ), .A1(\add_x_19_5/n116 ), .B0(
        \add_x_19_5/n117 ), .Y(\add_x_19_5/n115 ) );
  AOI21X4TS U1607 ( .A0(\add_x_19_5/n157 ), .A1(\add_x_19_5/n114 ), .B0(
        \add_x_19_5/n115 ), .Y(\add_x_19_5/n113 ) );
  OAI21X2TS U1608 ( .A0(\add_x_19_5/n113 ), .A1(\add_x_19_5/n93 ), .B0(
        \add_x_19_5/n94 ), .Y(\add_x_19_5/n92 ) );
  NOR2X4TS U1609 ( .A(n1883), .B(n2476), .Y(\add_x_19_3/n120 ) );
  NOR2X2TS U1610 ( .A(\add_x_19_3/n123 ), .B(\add_x_19_3/n120 ), .Y(
        \add_x_19_3/n118 ) );
  INVX1TS U1611 ( .A(\add_x_19_0/n73 ), .Y(\add_x_19_0/n71 ) );
  OAI21X2TS U1612 ( .A0(\add_x_19_0/n113 ), .A1(\add_x_19_0/n70 ), .B0(
        \add_x_19_0/n71 ), .Y(\add_x_19_0/n69 ) );
  INVX1TS U1613 ( .A(\add_x_19_0/n55 ), .Y(\add_x_19_0/n196 ) );
  NOR2X2TS U1614 ( .A(\add_x_19_4/n123 ), .B(\add_x_19_4/n120 ), .Y(n1549) );
  NAND2X2TS U1615 ( .A(\add_x_19_4/n126 ), .B(n1549), .Y(n1567) );
  NOR2X2TS U1616 ( .A(\addr_calc/fft_write_calc/count[5] ), .B(n2485), .Y(
        \add_x_19_1/n170 ) );
  NOR2X1TS U1617 ( .A(\add_x_19_3/n128 ), .B(\add_x_19_3/n131 ), .Y(
        \add_x_19_3/n126 ) );
  NOR2X2TS U1618 ( .A(n1990), .B(n2446), .Y(\add_x_19_3/n184 ) );
  AOI21X2TS U1619 ( .A0(\add_x_19_3/n179 ), .A1(\add_x_19_3/n187 ), .B0(
        \add_x_19_3/n180 ), .Y(\add_x_19_3/n178 ) );
  NOR2X2TS U1620 ( .A(n1967), .B(n2418), .Y(\add_x_19_0/n128 ) );
  NAND2X1TS U1621 ( .A(\add_x_19_3/n118 ), .B(\add_x_19_3/n126 ), .Y(
        \add_x_19_3/n116 ) );
  AOI2BB1X2TS U1622 ( .A0N(\add_x_19_1/n38 ), .A1N(n1550), .B0(n1551), .Y(
        \addr_calc/fft_write_addr[31] ) );
  OAI21X2TS U1623 ( .A0(\add_x_19_0/n191 ), .A1(\add_x_19_0/n188 ), .B0(
        \add_x_19_0/n189 ), .Y(\add_x_19_0/n187 ) );
  AOI21X2TS U1624 ( .A0(\add_x_19_1/n179 ), .A1(\add_x_19_1/n187 ), .B0(
        \add_x_19_1/n180 ), .Y(\add_x_19_1/n178 ) );
  INVX1TS U1625 ( .A(\add_x_19_1/n73 ), .Y(\add_x_19_1/n71 ) );
  INVX1TS U1626 ( .A(\add_x_19_1/n72 ), .Y(\add_x_19_1/n70 ) );
  AOI21X2TS U1627 ( .A0(\add_x_19_5/n112 ), .A1(\add_x_19_5/n103 ), .B0(
        \add_x_19_5/n104 ), .Y(\add_x_19_5/n102 ) );
  INVX1TS U1628 ( .A(\add_x_19_1/n55 ), .Y(\add_x_19_1/n196 ) );
  INVX1TS U1629 ( .A(\add_x_19_5/n97 ), .Y(\add_x_19_5/n204 ) );
  AOI21X1TS U1630 ( .A0(\add_x_19_0/n169 ), .A1(n1558), .B0(\add_x_19_0/n161 ), 
        .Y(\add_x_19_0/n159 ) );
  NAND2X1TS U1631 ( .A(n1558), .B(\add_x_19_0/n168 ), .Y(\add_x_19_0/n158 ) );
  AOI21X4TS U1632 ( .A0(\add_x_19_0/n157 ), .A1(\add_x_19_0/n114 ), .B0(
        \add_x_19_0/n115 ), .Y(\add_x_19_0/n113 ) );
  INVX2TS U1633 ( .A(\add_x_19_0/n157 ), .Y(\add_x_19_0/n156 ) );
  OAI21X2TS U1634 ( .A0(n1139), .A1(\add_x_19_0/n44 ), .B0(\add_x_19_0/n45 ), 
        .Y(\add_x_19_0/n43 ) );
  INVX2TS U1635 ( .A(\add_x_19_0/n113 ), .Y(\add_x_19_0/n112 ) );
  INVX1TS U1636 ( .A(\add_x_19_0/n92 ), .Y(\add_x_19_0/n91 ) );
  OAI21X1TS U1637 ( .A0(\add_x_19_0/n83 ), .A1(\add_x_19_0/n81 ), .B0(
        \add_x_19_0/n82 ), .Y(\add_x_19_0/n80 ) );
  XOR2X2TS U1638 ( .A(\add_x_19_0/n80 ), .B(n1561), .Y(
        \addr_calc/fft_read_addr[23] ) );
  OR2X1TS U1639 ( .A(\addr_calc/fir_read_calc/count[31] ), .B(n2380), .Y(n1560) );
  INVX1TS U1640 ( .A(\add_x_19_0/n78 ), .Y(\add_x_19_0/n200 ) );
  AND2X2TS U1641 ( .A(\add_x_19_0/n200 ), .B(\add_x_19_0/n79 ), .Y(n1561) );
  NOR2X2TS U1642 ( .A(\addr_calc/fir_write_calc/count[7] ), .B(n2422), .Y(
        \add_x_19_3/n162 ) );
  CLKINVX1TS U1643 ( .A(n2370), .Y(n1562) );
  INVX1TS U1644 ( .A(\DP_OP_159_297_3515/n902 ), .Y(\DP_OP_159_297_3515/n901 )
         );
  NAND2X2TS U1645 ( .A(n1791), .B(\DP_OP_159_297_3515/n900 ), .Y(
        \DP_OP_159_297_3515/n899 ) );
  XOR2X4TS U1646 ( .A(\DP_OP_159_297_3515/n899 ), .B(n1809), .Y(n2613) );
  XNOR2X4TS U1647 ( .A(n1738), .B(n2051), .Y(\DP_OP_159_297_3515/n541 ) );
  XNOR2X4TS U1648 ( .A(n1703), .B(n2579), .Y(\DP_OP_159_297_3515/n569 ) );
  XOR2X4TS U1649 ( .A(n1699), .B(n1961), .Y(\DP_OP_159_297_3515/n582 ) );
  XOR2X4TS U1650 ( .A(\DP_OP_159_297_3515/n1138 ), .B(
        \addr_calc/iir_write_calc/count[28] ), .Y(\DP_OP_159_297_3515/n476 )
         );
  XOR2X4TS U1651 ( .A(n1732), .B(n1968), .Y(\DP_OP_159_297_3515/n527 ) );
  XNOR2X4TS U1652 ( .A(n1661), .B(n2573), .Y(\DP_OP_159_297_3515/n512 ) );
  NOR2X4TS U1653 ( .A(\DP_OP_159_297_3515/n556 ), .B(\DP_OP_159_297_3515/n541 ), .Y(\DP_OP_159_297_3515/n539 ) );
  NOR2X4TS U1654 ( .A(\DP_OP_159_297_3515/n582 ), .B(\DP_OP_159_297_3515/n569 ), .Y(\DP_OP_159_297_3515/n567 ) );
  NOR2X4TS U1655 ( .A(\DP_OP_159_297_3515/n495 ), .B(\DP_OP_159_297_3515/n476 ), .Y(\DP_OP_159_297_3515/n474 ) );
  NOR2X4TS U1656 ( .A(\DP_OP_159_297_3515/n512 ), .B(\DP_OP_159_297_3515/n527 ), .Y(\DP_OP_159_297_3515/n510 ) );
  NAND2X2TS U1657 ( .A(n1564), .B(n1563), .Y(\DP_OP_159_297_3515/n443 ) );
  NAND2X4TS U1658 ( .A(\DP_OP_159_297_3515/n567 ), .B(
        \DP_OP_159_297_3515/n539 ), .Y(\DP_OP_159_297_3515/n537 ) );
  NAND2X4TS U1659 ( .A(\DP_OP_159_297_3515/n510 ), .B(
        \DP_OP_159_297_3515/n474 ), .Y(\DP_OP_159_297_3515/n472 ) );
  NOR2X2TS U1660 ( .A(\DP_OP_159_297_3515/n443 ), .B(\DP_OP_159_297_3515/n430 ), .Y(\DP_OP_159_297_3515/n428 ) );
  NOR2X4TS U1661 ( .A(\DP_OP_159_297_3515/n472 ), .B(\DP_OP_159_297_3515/n537 ), .Y(\DP_OP_159_297_3515/n470 ) );
  AND2X8TS U1662 ( .A(\DP_OP_159_297_3515/n470 ), .B(\DP_OP_159_297_3515/n428 ), .Y(n1779) );
  AOI21X4TS U1663 ( .A0(\addr_calc/iir_write_calc/counter/N38 ), .A1(
        data_from_iir), .B0(n1861), .Y(n2812) );
  OAI2BB1X2TS U1664 ( .A0N(n1951), .A1N(n2675), .B0(n1565), .Y(n986) );
  OAI21X2TS U1665 ( .A0(n1567), .A1(\add_x_19_4/n136 ), .B0(\add_x_19_4/n117 ), 
        .Y(\add_x_19_4/n115 ) );
  NOR2X2TS U1666 ( .A(n1567), .B(\add_x_19_4/n135 ), .Y(\add_x_19_4/n114 ) );
  AOI21X4TS U1667 ( .A0(\add_x_19_4/n157 ), .A1(\add_x_19_4/n114 ), .B0(
        \add_x_19_4/n115 ), .Y(\add_x_19_4/n113 ) );
  OAI21X2TS U1668 ( .A0(\add_x_19_4/n113 ), .A1(\add_x_19_4/n93 ), .B0(
        \add_x_19_4/n94 ), .Y(\add_x_19_4/n92 ) );
  OAI21X2TS U1669 ( .A0(\add_x_19_4/n113 ), .A1(\add_x_19_4/n44 ), .B0(
        \add_x_19_4/n45 ), .Y(\add_x_19_4/n43 ) );
  OAI21X2TS U1670 ( .A0(\add_x_19_4/n113 ), .A1(\add_x_19_4/n70 ), .B0(
        \add_x_19_4/n71 ), .Y(\add_x_19_4/n69 ) );
  INVX2TS U1671 ( .A(\add_x_19_4/n113 ), .Y(\add_x_19_4/n112 ) );
  AOI21X2TS U1672 ( .A0(\add_x_19_4/n92 ), .A1(\add_x_19_4/n84 ), .B0(
        \add_x_19_4/n85 ), .Y(\add_x_19_4/n83 ) );
  OAI21X2TS U1673 ( .A0(\add_x_19_4/n83 ), .A1(\add_x_19_4/n81 ), .B0(
        \add_x_19_4/n82 ), .Y(\add_x_19_4/n80 ) );
  OAI21X1TS U1674 ( .A0(\add_x_19_3/n155 ), .A1(\add_x_19_3/n151 ), .B0(
        \add_x_19_3/n152 ), .Y(\add_x_19_3/n150 ) );
  CLKINVX1TS U1675 ( .A(\add_x_19_4/n78 ), .Y(\add_x_19_4/n200 ) );
  XOR2X4TS U1676 ( .A(\add_x_19_4/n80 ), .B(n1466), .Y(
        \addr_calc/iir_read_addr[23] ) );
  OAI21X2TS U1677 ( .A0(\add_x_19_2/n91 ), .A1(\add_x_19_2/n89 ), .B0(
        \add_x_19_2/n90 ), .Y(n1568) );
  NAND2BX1TS U1678 ( .AN(n1571), .B(n1707), .Y(n1570) );
  OAI2BB1X1TS U1679 ( .A0N(n2576), .A1N(n2652), .B0(n1570), .Y(n945) );
  INVX1TS U1680 ( .A(\add_x_19_5/n78 ), .Y(\add_x_19_5/n200 ) );
  XNOR2X2TS U1681 ( .A(\add_x_19_5/n80 ), .B(\add_x_19_5/n9 ), .Y(
        \addr_calc/iir_write_addr[23] ) );
  OAI21X2TS U1682 ( .A0(\add_x_19_3/n132 ), .A1(\add_x_19_3/n128 ), .B0(
        \add_x_19_3/n129 ), .Y(\add_x_19_3/n127 ) );
  NAND2BX1TS U1683 ( .AN(n1574), .B(n1771), .Y(n1573) );
  OAI2BB1X2TS U1684 ( .A0N(n1948), .A1N(n2675), .B0(n1573), .Y(n987) );
  NAND2BX1TS U1685 ( .AN(n1577), .B(n1708), .Y(n1576) );
  OAI2BB1X1TS U1686 ( .A0N(n1929), .A1N(n2653), .B0(n1576), .Y(n944) );
  OAI21X1TS U1687 ( .A0(\add_x_19_4/n43 ), .A1(n1579), .B0(n1580), .Y(
        \addr_calc/iir_read_addr[30] ) );
  NOR2BX1TS U1688 ( .AN(n2634), .B(n1640), .Y(n1581) );
  AOI21X1TS U1689 ( .A0(\add_x_19_4/n43 ), .A1(n1581), .B0(n1582), .Y(n1580)
         );
  NAND2X1TS U1690 ( .A(n1640), .B(n1583), .Y(n1579) );
  OR2X2TS U1691 ( .A(n1847), .B(n2382), .Y(n1586) );
  NOR2XLTS U1692 ( .A(\add_x_19_0/n181 ), .B(\add_x_19_0/n184 ), .Y(n1587) );
  AOI21X1TS U1693 ( .A0(\add_x_19_0/n187 ), .A1(n1587), .B0(n1588), .Y(
        \add_x_19_0/n178 ) );
  OR2X2TS U1694 ( .A(\addr_calc/iir_write_calc/count[31] ), .B(n2381), .Y(
        n1590) );
  NOR2X1TS U1695 ( .A(\add_x_19_3/n135 ), .B(\add_x_19_3/n116 ), .Y(n1592) );
  AOI21X2TS U1696 ( .A0(\add_x_19_3/n157 ), .A1(n1592), .B0(n1593), .Y(
        \add_x_19_3/n113 ) );
  OAI21X1TS U1697 ( .A0(\add_x_19_3/n136 ), .A1(\add_x_19_3/n116 ), .B0(n1594), 
        .Y(n1593) );
  AOI21X2TS U1698 ( .A0(\add_x_19_3/n127 ), .A1(\add_x_19_3/n118 ), .B0(n1595), 
        .Y(n1594) );
  CLKINVX1TS U1699 ( .A(\add_x_19_3/n78 ), .Y(\add_x_19_3/n200 ) );
  OAI21X1TS U1700 ( .A0(\add_x_19_3/n83 ), .A1(\add_x_19_3/n81 ), .B0(
        \add_x_19_3/n82 ), .Y(\add_x_19_3/n80 ) );
  AOI21X2TS U1701 ( .A0(\add_x_19_2/n92 ), .A1(\add_x_19_2/n84 ), .B0(
        \add_x_19_2/n85 ), .Y(\add_x_19_2/n83 ) );
  NOR2X1TS U1702 ( .A(n1817), .B(n1508), .Y(\DP_OP_158_296_6262/n1850 ) );
  NAND2X2TS U1703 ( .A(\DP_OP_158_296_6262/n1862 ), .B(
        \DP_OP_158_296_6262/n1850 ), .Y(\DP_OP_158_296_6262/n1792 ) );
  XOR2X1TS U1704 ( .A(n2596), .B(\addr_calc/fft_read_calc/count[2] ), .Y(n1598) );
  XOR2X1TS U1705 ( .A(\DP_OP_158_296_6262/n855 ), .B(
        \addr_calc/fft_read_calc/count[4] ), .Y(n1601) );
  XOR2X1TS U1706 ( .A(n2599), .B(n1978), .Y(n1600) );
  XOR2X1TS U1707 ( .A(n2593), .B(\addr_calc/fft_read_calc/count[6] ), .Y(n1599) );
  XNOR2X2TS U1708 ( .A(n1660), .B(n1970), .Y(\DP_OP_158_296_6262/n1180 ) );
  XOR2X4TS U1709 ( .A(n1654), .B(n1955), .Y(\DP_OP_158_296_6262/n1079 ) );
  XNOR2X1TS U1710 ( .A(n1775), .B(\addr_calc/fft_read_calc/count[28] ), .Y(
        \DP_OP_158_296_6262/n948 ) );
  XOR2X4TS U1711 ( .A(n1718), .B(n2037), .Y(\DP_OP_158_296_6262/n1013 ) );
  XOR2X4TS U1712 ( .A(\DP_OP_158_296_6262/n833 ), .B(\add_x_22_0/n15 ), .Y(
        \DP_OP_158_296_6262/n981 ) );
  XNOR2X2TS U1713 ( .A(n1776), .B(n2572), .Y(\DP_OP_158_296_6262/n1068 ) );
  NOR2X2TS U1714 ( .A(\DP_OP_158_296_6262/n1243 ), .B(
        \DP_OP_158_296_6262/n1259 ), .Y(\DP_OP_158_296_6262/n1241 ) );
  NOR2X2TS U1715 ( .A(\DP_OP_158_296_6262/n1216 ), .B(
        \DP_OP_158_296_6262/n1223 ), .Y(\DP_OP_158_296_6262/n1214 ) );
  NOR2X2TS U1716 ( .A(\DP_OP_158_296_6262/n1200 ), .B(
        \DP_OP_158_296_6262/n1209 ), .Y(\DP_OP_158_296_6262/n1198 ) );
  NOR2X2TS U1717 ( .A(\DP_OP_158_296_6262/n1191 ), .B(
        \DP_OP_158_296_6262/n1180 ), .Y(\DP_OP_158_296_6262/n1178 ) );
  NOR2X2TS U1718 ( .A(\DP_OP_158_296_6262/n1149 ), .B(
        \DP_OP_158_296_6262/n1136 ), .Y(\DP_OP_158_296_6262/n1134 ) );
  NOR2X2TS U1719 ( .A(\DP_OP_158_296_6262/n933 ), .B(\DP_OP_158_296_6262/n948 ), .Y(\DP_OP_158_296_6262/n931 ) );
  NOR2X4TS U1720 ( .A(\DP_OP_158_296_6262/n981 ), .B(\DP_OP_158_296_6262/n962 ), .Y(\DP_OP_158_296_6262/n960 ) );
  NOR2X4TS U1721 ( .A(\DP_OP_158_296_6262/n1042 ), .B(
        \DP_OP_158_296_6262/n1027 ), .Y(\DP_OP_158_296_6262/n1025 ) );
  NOR2X4TS U1722 ( .A(\DP_OP_158_296_6262/n1068 ), .B(
        \DP_OP_158_296_6262/n1055 ), .Y(\DP_OP_158_296_6262/n1053 ) );
  NAND2X2TS U1723 ( .A(\DP_OP_158_296_6262/n1214 ), .B(
        \DP_OP_158_296_6262/n1241 ), .Y(\DP_OP_158_296_6262/n1212 ) );
  NAND2X2TS U1724 ( .A(\DP_OP_158_296_6262/n1178 ), .B(
        \DP_OP_158_296_6262/n1198 ), .Y(\DP_OP_158_296_6262/n1176 ) );
  NAND2X2TS U1725 ( .A(\DP_OP_158_296_6262/n1158 ), .B(
        \DP_OP_158_296_6262/n1134 ), .Y(\DP_OP_158_296_6262/n1132 ) );
  NAND2X2TS U1726 ( .A(\DP_OP_158_296_6262/n1077 ), .B(
        \DP_OP_158_296_6262/n1109 ), .Y(\DP_OP_158_296_6262/n1075 ) );
  NAND2X2TS U1727 ( .A(\DP_OP_158_296_6262/n931 ), .B(n1471), .Y(
        \DP_OP_158_296_6262/n912 ) );
  NOR2X2TS U1728 ( .A(\DP_OP_158_296_6262/n912 ), .B(\DP_OP_158_296_6262/n899 ), .Y(\DP_OP_158_296_6262/n897 ) );
  NAND2X2TS U1729 ( .A(\DP_OP_158_296_6262/n897 ), .B(
        \DP_OP_158_296_6262/n956 ), .Y(\DP_OP_158_296_6262/n895 ) );
  OR2X8TS U1730 ( .A(\DP_OP_158_296_6262/n895 ), .B(\DP_OP_158_296_6262/n1071 ), .Y(\addr_calc/fft_read_calc/counter/N38 ) );
  AOI21X4TS U1731 ( .A0(\addr_calc/fft_read_calc/counter/N38 ), .A1(
        data_to_fft), .B0(n2588), .Y(n2794) );
  OAI2BB1X2TS U1732 ( .A0N(n1605), .A1N(\add_x_19_5/n60 ), .B0(n1606), .Y(
        n1604) );
  AOI2BB1X2TS U1733 ( .A0N(\add_x_19_5/n60 ), .A1N(n1603), .B0(n1604), .Y(
        \addr_calc/iir_write_addr[27] ) );
  NAND2BX1TS U1734 ( .AN(n1609), .B(n1751), .Y(n1608) );
  NOR2X4TS U1735 ( .A(n1813), .B(n1529), .Y(\DP_OP_158_296_6262/n1918 ) );
  INVX2TS U1736 ( .A(\add_x_19_4/n69 ), .Y(n1611) );
  XNOR2X1TS U1737 ( .A(n1611), .B(n1467), .Y(\addr_calc/iir_read_addr[24] ) );
  OAI21X2TS U1738 ( .A0(n1611), .A1(\add_x_19_4/n51 ), .B0(\add_x_19_4/n52 ), 
        .Y(\add_x_19_4/n50 ) );
  OAI21X2TS U1739 ( .A0(n1611), .A1(\add_x_19_4/n66 ), .B0(\add_x_19_4/n67 ), 
        .Y(\add_x_19_4/n65 ) );
  NAND2X4TS U1740 ( .A(\DP_OP_158_296_6262/n1918 ), .B(
        \DP_OP_158_296_6262/n1906 ), .Y(\DP_OP_158_296_6262/n1903 ) );
  INVXLTS U1741 ( .A(\DP_OP_158_296_6262/n1890 ), .Y(
        \DP_OP_158_296_6262/n1891 ) );
  XNOR2X4TS U1742 ( .A(\DP_OP_158_296_6262/n1881 ), .B(n2344), .Y(n1730) );
  AOI21X4TS U1743 ( .A0(\addr_calc/fir_write_calc/counter/N38 ), .A1(
        data_from_fir), .B0(n2061), .Y(n2805) );
  NAND2BX1TS U1744 ( .AN(n1613), .B(n1826), .Y(n1612) );
  NAND2X1TS U1745 ( .A(n1763), .B(\addr_calc/fir_write_calc/counter/N73 ), .Y(
        n1617) );
  OAI2BB1X1TS U1746 ( .A0N(n1836), .A1N(n1262), .B0(n1617), .Y(n1100) );
  NAND2BX1TS U1747 ( .AN(n1619), .B(n1764), .Y(n1618) );
  OAI2BB1X2TS U1748 ( .A0N(n1970), .A1N(n2657), .B0(n1620), .Y(n1023) );
  INVX2TS U1749 ( .A(n2344), .Y(\DP_OP_159_297_3515/n861 ) );
  NAND2X2TS U1750 ( .A(n1790), .B(\DP_OP_159_297_3515/n942 ), .Y(
        \DP_OP_159_297_3515/n941 ) );
  XOR2X4TS U1751 ( .A(\DP_OP_159_297_3515/n941 ), .B(\DP_OP_159_297_3515/n861 ), .Y(\DP_OP_159_297_3515/n1133 ) );
  XOR2X4TS U1752 ( .A(n1703), .B(\add_x_22_4/n33 ), .Y(
        \DP_OP_159_297_3515/n144 ) );
  XOR2X4TS U1753 ( .A(n1699), .B(n1923), .Y(\DP_OP_159_297_3515/n157 ) );
  XOR2X4TS U1754 ( .A(\DP_OP_159_297_3515/n1138 ), .B(
        \addr_calc/iir_read_calc/count[28] ), .Y(\DP_OP_159_297_3515/n51 ) );
  XNOR2X4TS U1755 ( .A(n1702), .B(\addr_calc/iir_read_calc/count[27] ), .Y(
        \DP_OP_159_297_3515/n70 ) );
  XOR2X4TS U1756 ( .A(n1732), .B(n1925), .Y(\DP_OP_159_297_3515/n102 ) );
  NOR2X4TS U1757 ( .A(\DP_OP_159_297_3515/n131 ), .B(\DP_OP_159_297_3515/n116 ), .Y(\DP_OP_159_297_3515/n114 ) );
  NOR2X4TS U1758 ( .A(\DP_OP_159_297_3515/n144 ), .B(\DP_OP_159_297_3515/n157 ), .Y(\DP_OP_159_297_3515/n142 ) );
  NOR2X4TS U1759 ( .A(\DP_OP_159_297_3515/n70 ), .B(\DP_OP_159_297_3515/n51 ), 
        .Y(\DP_OP_159_297_3515/n49 ) );
  NAND2X4TS U1760 ( .A(\DP_OP_159_297_3515/n114 ), .B(
        \DP_OP_159_297_3515/n142 ), .Y(\DP_OP_159_297_3515/n112 ) );
  NAND2X4TS U1761 ( .A(\DP_OP_159_297_3515/n85 ), .B(\DP_OP_159_297_3515/n49 ), 
        .Y(\DP_OP_159_297_3515/n47 ) );
  NOR2X4TS U1762 ( .A(\DP_OP_159_297_3515/n18 ), .B(\DP_OP_159_297_3515/n5 ), 
        .Y(\DP_OP_159_297_3515/n3 ) );
  NOR2X8TS U1763 ( .A(\DP_OP_159_297_3515/n47 ), .B(\DP_OP_159_297_3515/n112 ), 
        .Y(\DP_OP_159_297_3515/n45 ) );
  NAND2X4TS U1764 ( .A(\DP_OP_159_297_3515/n45 ), .B(\DP_OP_159_297_3515/n3 ), 
        .Y(\DP_OP_159_297_3515/n1 ) );
  NOR2BX4TS U1765 ( .AN(n1625), .B(n1675), .Y(n2795) );
  OAI2BB1X2TS U1766 ( .A0N(n1953), .A1N(n1476), .B0(n1627), .Y(n1013) );
  NAND2BX1TS U1767 ( .AN(n1631), .B(n1754), .Y(n1630) );
  OAI2BB1X2TS U1768 ( .A0N(n2575), .A1N(n1477), .B0(n1630), .Y(n1008) );
  INVX2TS U1769 ( .A(\add_x_19_4/n128 ), .Y(n1632) );
  NAND2BX1TS U1770 ( .AN(n1634), .B(n1751), .Y(n1633) );
  OAI2BB1X2TS U1771 ( .A0N(\addr_calc/fft_read_calc/count[17] ), .A1N(n1475), 
        .B0(n1633), .Y(n1017) );
  NOR2X4TS U1772 ( .A(filesize[1]), .B(n1525), .Y(n1797) );
  OAI21X2TS U1773 ( .A0(\add_x_19_4/n156 ), .A1(\add_x_19_4/n135 ), .B0(
        \add_x_19_4/n136 ), .Y(\add_x_19_4/n134 ) );
  CLKINVX1TS U1774 ( .A(\add_x_19_4/n120 ), .Y(\add_x_19_4/n208 ) );
  NAND2BX1TS U1775 ( .AN(n1637), .B(n1754), .Y(n1636) );
  OAI2BB1X2TS U1776 ( .A0N(n2569), .A1N(n1476), .B0(n1636), .Y(n1016) );
  NAND2BX1TS U1777 ( .AN(n1639), .B(n1749), .Y(n1638) );
  OAI2BB1X2TS U1778 ( .A0N(n2554), .A1N(n1475), .B0(n1638), .Y(n1018) );
  AOI21X1TS U1779 ( .A0(\add_x_19_4/n73 ), .A1(\add_x_19_4/n46 ), .B0(
        \add_x_19_4/n47 ), .Y(\add_x_19_4/n45 ) );
  INVX2TS U1780 ( .A(\add_x_19_4/n42 ), .Y(\add_x_19_4/n40 ) );
  CLKINVX2TS U1781 ( .A(\add_x_19_4/n72 ), .Y(\add_x_19_4/n70 ) );
  INVX1TS U1782 ( .A(\add_x_19_4/n63 ), .Y(\add_x_19_4/n198 ) );
  CLKINVX1TS U1783 ( .A(\add_x_19_4/n48 ), .Y(\add_x_19_4/n195 ) );
  XOR2X4TS U1784 ( .A(\DP_OP_158_296_6262/n1860 ), .B(n1664), .Y(
        \DP_OP_158_296_6262/n2056 ) );
  XOR2X4TS U1785 ( .A(n1642), .B(\DP_OP_158_296_6262/n1897 ), .Y(n1776) );
  NAND2BX1TS U1786 ( .AN(n1644), .B(n1751), .Y(n1643) );
  OAI2BB1X2TS U1787 ( .A0N(n2552), .A1N(n2656), .B0(n1643), .Y(n1030) );
  NAND2BX1TS U1788 ( .AN(n1837), .B(n1744), .Y(n1645) );
  NAND2BX1TS U1789 ( .AN(n1647), .B(n1763), .Y(n1646) );
  OAI2BB1X2TS U1790 ( .A0N(n2000), .A1N(n1264), .B0(n1646), .Y(n1118) );
  NOR2X2TS U1791 ( .A(filesize[1]), .B(filesize[2]), .Y(
        \DP_OP_159_297_3515/n1075 ) );
  NAND2X1TS U1792 ( .A(n1527), .B(n1497), .Y(\DP_OP_159_297_3515/n1066 ) );
  XOR2X2TS U1793 ( .A(n1790), .B(\DP_OP_159_297_3515/n867 ), .Y(n2607) );
  CLKBUFX2TS U1794 ( .A(n1525), .Y(n1648) );
  AO22X4TS U1795 ( .A0(n1773), .A1(\addr_calc/iir_write_calc/counter/N60 ), 
        .B0(n1954), .B1(n2676), .Y(n985) );
  BUFX6TS U1796 ( .A(n2679), .Y(n2676) );
  AO22X4TS U1797 ( .A0(n1772), .A1(\addr_calc/iir_write_calc/counter/N66 ), 
        .B0(n2674), .B1(\addr_calc/iir_write_calc/count[23] ), .Y(n979) );
  AO22X4TS U1798 ( .A0(n1769), .A1(\addr_calc/iir_write_calc/counter/N74 ), 
        .B0(n2675), .B1(n1857), .Y(n1136) );
  XNOR2X2TS U1799 ( .A(\add_x_19_4/n88 ), .B(\add_x_19_4/n11 ), .Y(
        \addr_calc/iir_read_addr[21] ) );
  BUFX8TS U1800 ( .A(n2679), .Y(n2672) );
  AO22X4TS U1801 ( .A0(n1770), .A1(\addr_calc/iir_write_calc/counter/N44 ), 
        .B0(n2677), .B1(n1931), .Y(n1001) );
  AO22X4TS U1802 ( .A0(n1771), .A1(\addr_calc/iir_write_calc/counter/N67 ), 
        .B0(n2677), .B1(\addr_calc/iir_write_calc/count[24] ), .Y(n978) );
  AO22X4TS U1803 ( .A0(n1772), .A1(\addr_calc/iir_write_calc/counter/N46 ), 
        .B0(n2677), .B1(n1933), .Y(n999) );
  AO22X4TS U1804 ( .A0(n1768), .A1(\addr_calc/iir_write_calc/counter/N48 ), 
        .B0(n2677), .B1(n1686), .Y(n997) );
  NOR2X6TS U1805 ( .A(n1468), .B(n787), .Y(n2813) );
  NOR2X1TS U1806 ( .A(n2789), .B(n2788), .Y(n2790) );
  INVX8TS U1807 ( .A(n2673), .Y(n1740) );
  OAI2BB2X2TS U1808 ( .B0(n1740), .B1(\add_x_22_5/n117 ), .A0N(n1773), .A1N(
        \addr_calc/iir_write_calc/counter/N45 ), .Y(n1000) );
  NAND2X2TS U1809 ( .A(n1792), .B(\DP_OP_159_297_3515/n928 ), .Y(
        \DP_OP_159_297_3515/n927 ) );
  NAND2X2TS U1810 ( .A(n1792), .B(\DP_OP_159_297_3515/n956 ), .Y(
        \DP_OP_159_297_3515/n955 ) );
  BUFX6TS U1811 ( .A(n2680), .Y(n2674) );
  NAND2X4TS U1812 ( .A(n1779), .B(n1780), .Y(n1649) );
  XOR2X4TS U1813 ( .A(\DP_OP_159_297_3515/n927 ), .B(n1484), .Y(n1732) );
  OAI2BB2X4TS U1814 ( .B0(n1740), .B1(n1973), .A0N(n1767), .A1N(
        \addr_calc/iir_write_calc/counter/N71 ), .Y(n974) );
  NOR4XLTS U1815 ( .A(n1478), .B(iir_write_done), .C(n925), .D(n926), .Y(n796)
         );
  AO22X4TS U1816 ( .A0(n1774), .A1(\addr_calc/iir_write_calc/counter/N49 ), 
        .B0(n2673), .B1(n2039), .Y(n996) );
  NOR2X4TS U1817 ( .A(\DP_OP_158_296_6262/n1903 ), .B(
        \DP_OP_158_296_6262/n1877 ), .Y(n1783) );
  XNOR2X1TS U1818 ( .A(n1776), .B(n1985), .Y(\DP_OP_158_296_6262/n174 ) );
  NOR2XLTS U1819 ( .A(filesize[1]), .B(filesize[2]), .Y(n1650) );
  XNOR2X4TS U1820 ( .A(\DP_OP_158_296_6262/n1991 ), .B(n2362), .Y(n1651) );
  XNOR2X4TS U1821 ( .A(\DP_OP_158_296_6262/n1909 ), .B(n1531), .Y(n1654) );
  XNOR2X4TS U1822 ( .A(\DP_OP_158_296_6262/n1971 ), .B(n2367), .Y(n1656) );
  XNOR2X4TS U1823 ( .A(\DP_OP_158_296_6262/n1943 ), .B(n1831), .Y(n1657) );
  XNOR2X4TS U1824 ( .A(\DP_OP_158_296_6262/n1936 ), .B(n1521), .Y(n1658) );
  XNOR2X4TS U1825 ( .A(\DP_OP_158_296_6262/n1964 ), .B(n1681), .Y(n1660) );
  XNOR2X4TS U1826 ( .A(\DP_OP_159_297_3515/n920 ), .B(n2343), .Y(n1661) );
  AOI21X2TS U1827 ( .A0(\add_x_19_4/n112 ), .A1(\add_x_19_4/n103 ), .B0(
        \add_x_19_4/n104 ), .Y(\add_x_19_4/n102 ) );
  BUFX8TS U1828 ( .A(n2679), .Y(n2678) );
  BUFX8TS U1829 ( .A(n2680), .Y(n2677) );
  NAND2X2TS U1830 ( .A(n1788), .B(\DP_OP_159_297_3515/n1011 ), .Y(
        \DP_OP_159_297_3515/n1010 ) );
  XNOR2X4TS U1831 ( .A(\DP_OP_159_297_3515/n1003 ), .B(
        \DP_OP_159_297_3515/n870 ), .Y(n2617) );
  XOR2X2TS U1832 ( .A(\DP_OP_158_296_6262/n2010 ), .B(n2371), .Y(
        \DP_OP_158_296_6262/n2034 ) );
  NOR2X4TS U1833 ( .A(n1717), .B(\DP_OP_158_296_6262/n1875 ), .Y(
        \DP_OP_158_296_6262/n1874 ) );
  NAND2X2TS U1834 ( .A(n1792), .B(\DP_OP_159_297_3515/n949 ), .Y(
        \DP_OP_159_297_3515/n948 ) );
  CLKINVX3TS U1835 ( .A(n1782), .Y(n1791) );
  INVX2TS U1836 ( .A(n1719), .Y(n1725) );
  INVX2TS U1837 ( .A(n1820), .Y(n1825) );
  INVX3TS U1838 ( .A(n1766), .Y(n1772) );
  INVX2TS U1839 ( .A(n1704), .Y(n1755) );
  INVX1TS U1840 ( .A(\add_x_19_2/n92 ), .Y(\add_x_19_2/n91 ) );
  CLKINVX2TS U1841 ( .A(\add_x_22_2/n24 ), .Y(\add_x_22_2/n23 ) );
  CLKINVX2TS U1842 ( .A(\add_x_22_5/n24 ), .Y(\add_x_22_5/n23 ) );
  CLKINVX2TS U1843 ( .A(\add_x_22_3/n24 ), .Y(\add_x_22_3/n23 ) );
  CLKINVX2TS U1844 ( .A(\add_x_22_5/n76 ), .Y(\add_x_22_5/n75 ) );
  INVX2TS U1845 ( .A(\add_x_22_4/n24 ), .Y(\add_x_22_4/n23 ) );
  CLKINVX2TS U1846 ( .A(\add_x_22_4/n42 ), .Y(\add_x_22_4/n41 ) );
  CLKINVX2TS U1847 ( .A(\add_x_22_3/n76 ), .Y(\add_x_22_3/n75 ) );
  INVX1TS U1848 ( .A(\add_x_22_4/n76 ), .Y(\add_x_22_4/n75 ) );
  CLKINVX2TS U1849 ( .A(\add_x_22_1/n24 ), .Y(\add_x_22_1/n23 ) );
  XNOR2X1TS U1850 ( .A(n1756), .B(n1994), .Y(\DP_OP_158_296_6262/n277 ) );
  INVX2TS U1851 ( .A(\add_x_22_0/n94 ), .Y(\add_x_22_0/n93 ) );
  NOR2X1TS U1852 ( .A(\add_x_19_4/n93 ), .B(\add_x_19_4/n74 ), .Y(
        \add_x_19_4/n72 ) );
  CLKINVX2TS U1853 ( .A(\add_x_19_3/n178 ), .Y(\add_x_19_3/n177 ) );
  NOR2X1TS U1854 ( .A(n2551), .B(n1155), .Y(\DP_OP_159_297_3515/n921 ) );
  CLKINVX1TS U1855 ( .A(\add_x_22_5/n119 ), .Y(\add_x_22_5/n118 ) );
  INVX1TS U1856 ( .A(\add_x_19_3/n176 ), .Y(\add_x_19_3/n174 ) );
  CLKINVX1TS U1857 ( .A(\add_x_19_4/n145 ), .Y(\add_x_19_4/n143 ) );
  INVX1TS U1858 ( .A(n1515), .Y(\DP_OP_159_297_3515/n862 ) );
  INVX1TS U1859 ( .A(\add_x_19_1/n144 ), .Y(\add_x_19_1/n213 ) );
  CLKINVX1TS U1860 ( .A(\add_x_19_1/n145 ), .Y(\add_x_19_1/n143 ) );
  CLKINVX1TS U1861 ( .A(\add_x_19_0/n175 ), .Y(\add_x_19_0/n219 ) );
  CLKINVX1TS U1862 ( .A(\add_x_19_3/n48 ), .Y(\add_x_19_3/n195 ) );
  CLKINVX1TS U1863 ( .A(\add_x_19_1/n48 ), .Y(\add_x_19_1/n195 ) );
  INVX1TS U1864 ( .A(\add_x_19_0/n48 ), .Y(\add_x_19_0/n195 ) );
  INVX2TS U1865 ( .A(n2013), .Y(n2014) );
  INVX2TS U1866 ( .A(n1901), .Y(n1902) );
  INVX2TS U1867 ( .A(n2045), .Y(n2046) );
  INVX2TS U1868 ( .A(n1975), .Y(n1666) );
  INVX2TS U1869 ( .A(\addr_calc/iir_read_calc/count[9] ), .Y(n1907) );
  INVX2TS U1870 ( .A(\addr_calc/iir_read_calc/count[18] ), .Y(n2024) );
  INVX2TS U1871 ( .A(\addr_calc/iir_write_calc/count[18] ), .Y(
        \add_x_22_5/n49 ) );
  INVX2TS U1872 ( .A(\addr_calc/iir_write_calc/count[14] ), .Y(
        \add_x_22_5/n67 ) );
  INVX2TS U1873 ( .A(\addr_calc/iir_read_calc/count[27] ), .Y(n1928) );
  INVX2TS U1874 ( .A(\addr_calc/fft_write_calc/count[19] ), .Y(n1921) );
  INVX2TS U1875 ( .A(\addr_calc/fir_write_calc/count[21] ), .Y(n1891) );
  INVX2TS U1876 ( .A(\addr_calc/fir_read_calc/count[22] ), .Y(n1981) );
  INVX2TS U1877 ( .A(\addr_calc/iir_write_calc/count[7] ), .Y(n1938) );
  BUFX3TS U1878 ( .A(\addr_calc/fir_write_calc/count[6] ), .Y(n1992) );
  BUFX3TS U1879 ( .A(\addr_calc/fir_write_calc/count[8] ), .Y(n1995) );
  INVX1TS U1880 ( .A(n2411), .Y(n2414) );
  INVX1TS U1881 ( .A(n2427), .Y(n2429) );
  INVX1TS U1882 ( .A(n2391), .Y(n2394) );
  CLKINVX1TS U1883 ( .A(n2391), .Y(n2393) );
  CLKINVX1TS U1884 ( .A(n2312), .Y(n2313) );
  INVX1TS U1885 ( .A(n2375), .Y(n2377) );
  INVX1TS U1886 ( .A(n2439), .Y(n2440) );
  INVX1TS U1887 ( .A(n2435), .Y(n2438) );
  INVX1TS U1888 ( .A(n2490), .Y(n2492) );
  INVX4TS U1889 ( .A(n1704), .Y(n1750) );
  INVX3TS U1890 ( .A(n1745), .Y(n1663) );
  INVX2TS U1891 ( .A(\add_x_19_3/n69 ), .Y(\add_x_19_3/n68 ) );
  NAND2X2TS U1892 ( .A(n1733), .B(n1681), .Y(n1735) );
  INVX1TS U1893 ( .A(\add_x_22_2/n76 ), .Y(\add_x_22_2/n75 ) );
  INVX1TS U1894 ( .A(\add_x_22_0/n76 ), .Y(\add_x_22_0/n75 ) );
  INVX1TS U1895 ( .A(\add_x_22_1/n76 ), .Y(\add_x_22_1/n75 ) );
  CLKINVX2TS U1896 ( .A(\add_x_19_3/n72 ), .Y(\add_x_19_3/n70 ) );
  NOR2X1TS U1897 ( .A(\add_x_19_3/n51 ), .B(\add_x_19_3/n48 ), .Y(
        \add_x_19_3/n46 ) );
  CLKINVX2TS U1898 ( .A(\add_x_19_5/n73 ), .Y(\add_x_19_5/n71 ) );
  OAI21X1TS U1899 ( .A0(\add_x_19_1/n94 ), .A1(\add_x_19_1/n74 ), .B0(
        \add_x_19_1/n75 ), .Y(\add_x_19_1/n73 ) );
  INVX1TS U1900 ( .A(\add_x_19_0/n178 ), .Y(\add_x_19_0/n177 ) );
  NAND2X1TS U1901 ( .A(\add_x_19_3/n61 ), .B(\add_x_19_3/n53 ), .Y(
        \add_x_19_3/n51 ) );
  NOR2X1TS U1902 ( .A(\add_x_19_3/n93 ), .B(\add_x_19_3/n74 ), .Y(
        \add_x_19_3/n72 ) );
  OAI21X1TS U1903 ( .A0(\add_x_19_4/n94 ), .A1(\add_x_19_4/n74 ), .B0(
        \add_x_19_4/n75 ), .Y(\add_x_19_4/n73 ) );
  INVX1TS U1904 ( .A(\add_x_19_2/n150 ), .Y(\add_x_19_2/n148 ) );
  INVX1TS U1905 ( .A(\add_x_19_1/n150 ), .Y(\add_x_19_1/n148 ) );
  INVX1TS U1906 ( .A(\add_x_19_3/n150 ), .Y(\add_x_19_3/n148 ) );
  INVX1TS U1907 ( .A(\add_x_19_0/n150 ), .Y(\add_x_19_0/n148 ) );
  INVX1TS U1908 ( .A(\add_x_19_2/n178 ), .Y(\add_x_19_2/n177 ) );
  INVX1TS U1909 ( .A(\add_x_19_0/n187 ), .Y(\add_x_19_0/n186 ) );
  INVX1TS U1910 ( .A(\add_x_19_5/n48 ), .Y(\add_x_19_5/n195 ) );
  CLKINVX1TS U1911 ( .A(\add_x_19_4/n55 ), .Y(\add_x_19_4/n196 ) );
  INVX2TS U1912 ( .A(n2066), .Y(n2061) );
  INVX1TS U1913 ( .A(\add_x_19_1/n187 ), .Y(\add_x_19_1/n186 ) );
  INVX1TS U1914 ( .A(\add_x_19_2/n111 ), .Y(\add_x_19_2/n109 ) );
  INVX1TS U1915 ( .A(\add_x_19_2/n187 ), .Y(\add_x_19_2/n186 ) );
  INVX1TS U1916 ( .A(\add_x_19_2/n144 ), .Y(\add_x_19_2/n213 ) );
  INVX1TS U1917 ( .A(\add_x_19_3/n187 ), .Y(\add_x_19_3/n186 ) );
  NOR2X1TS U1918 ( .A(\add_x_19_0/n58 ), .B(\add_x_19_0/n55 ), .Y(
        \add_x_19_0/n53 ) );
  NOR2X2TS U1919 ( .A(n1685), .B(n1980), .Y(\add_x_19_4/n151 ) );
  INVX1TS U1920 ( .A(\add_x_19_5/n187 ), .Y(\add_x_19_5/n186 ) );
  INVX1TS U1921 ( .A(\add_x_19_5/n175 ), .Y(\add_x_19_5/n219 ) );
  INVX1TS U1922 ( .A(\add_x_19_1/n111 ), .Y(\add_x_19_1/n109 ) );
  NOR2X1TS U1923 ( .A(\add_x_19_4/n81 ), .B(\add_x_19_4/n78 ), .Y(
        \add_x_19_4/n76 ) );
  NOR2X1TS U1924 ( .A(\add_x_19_5/n110 ), .B(\add_x_19_5/n105 ), .Y(
        \add_x_19_5/n103 ) );
  INVX1TS U1925 ( .A(\add_x_19_4/n188 ), .Y(\add_x_19_4/n222 ) );
  INVX1TS U1926 ( .A(\add_x_19_5/n188 ), .Y(\add_x_19_5/n222 ) );
  INVX1TS U1927 ( .A(\add_x_19_0/n144 ), .Y(\add_x_19_0/n213 ) );
  INVX1TS U1928 ( .A(\add_x_19_1/n175 ), .Y(\add_x_19_1/n219 ) );
  INVX1TS U1929 ( .A(\add_x_19_0/n111 ), .Y(\add_x_19_0/n109 ) );
  INVX1TS U1930 ( .A(\add_x_19_4/n175 ), .Y(\add_x_19_4/n219 ) );
  INVX2TS U1931 ( .A(\DP_OP_159_297_3515/n875 ), .Y(n2365) );
  INVX2TS U1932 ( .A(n801), .Y(n2053) );
  INVX2TS U1933 ( .A(\DP_OP_159_297_3515/n876 ), .Y(n2364) );
  INVX2TS U1934 ( .A(\DP_OP_159_297_3515/n868 ), .Y(n2361) );
  INVX2TS U1935 ( .A(\DP_OP_159_297_3515/n878 ), .Y(n2366) );
  INVX2TS U1936 ( .A(n1837), .Y(n1838) );
  INVX2TS U1937 ( .A(n2016), .Y(n2017) );
  INVX2TS U1938 ( .A(\add_x_22_4/n67 ), .Y(n1784) );
  INVX2TS U1939 ( .A(n1982), .Y(n1983) );
  INVX2TS U1940 ( .A(n1984), .Y(n1985) );
  INVX2TS U1941 ( .A(n1991), .Y(n1690) );
  INVX2TS U1942 ( .A(\add_x_22_4/n64 ), .Y(n2566) );
  INVX2TS U1943 ( .A(n1834), .Y(n1835) );
  INVX2TS U1944 ( .A(n1937), .Y(n1686) );
  INVX2TS U1945 ( .A(n1998), .Y(n2000) );
  INVX2TS U1946 ( .A(n2042), .Y(n2043) );
  INVX2TS U1947 ( .A(n1963), .Y(n1689) );
  INVX1TS U1948 ( .A(n1903), .Y(\add_x_22_4/n109 ) );
  CLKINVX2TS U1949 ( .A(n1955), .Y(n1956) );
  INVX2TS U1950 ( .A(\add_x_22_0/n49 ), .Y(n2569) );
  INVX2TS U1951 ( .A(n1850), .Y(n1851) );
  INVX2TS U1952 ( .A(n2027), .Y(n2028) );
  CLKINVX4TS U1953 ( .A(n2343), .Y(n1664) );
  NOR2X1TS U1954 ( .A(n1809), .B(n1807), .Y(\DP_OP_158_296_6262/n1837 ) );
  INVX2TS U1955 ( .A(\addr_calc/fft_write_calc/count[30] ), .Y(n1848) );
  INVX2TS U1956 ( .A(\addr_calc/fft_read_calc/count[3] ), .Y(\add_x_22_0/n114 ) );
  BUFX3TS U1957 ( .A(\addr_calc/iir_write_calc/count[3] ), .Y(n1933) );
  BUFX3TS U1958 ( .A(\addr_calc/fir_write_calc/count[4] ), .Y(n1865) );
  INVX2TS U1959 ( .A(\addr_calc/iir_write_calc/count[5] ), .Y(n1937) );
  INVX2TS U1960 ( .A(\addr_calc/fft_read_calc/count[30] ), .Y(n1858) );
  INVX2TS U1961 ( .A(\addr_calc/iir_write_calc/count[20] ), .Y(n2047) );
  INVX2TS U1962 ( .A(n2040), .Y(n1665) );
  INVX2TS U1963 ( .A(\addr_calc/fft_read_calc/count[21] ), .Y(n1952) );
  INVX2TS U1964 ( .A(\addr_calc/iir_read_calc/count[21] ), .Y(n1923) );
  INVX2TS U1965 ( .A(\addr_calc/iir_write_calc/count[27] ), .Y(n1971) );
  BUFX3TS U1966 ( .A(\addr_calc/iir_read_calc/count[11] ), .Y(n1911) );
  INVX2TS U1967 ( .A(\addr_calc/fft_read_calc/count[26] ), .Y(\add_x_22_0/n15 ) );
  BUFX3TS U1968 ( .A(\addr_calc/fft_write_calc/count[0] ), .Y(n2035) );
  INVX2TS U1969 ( .A(\addr_calc/iir_read_calc/count[19] ), .Y(\add_x_22_4/n46 ) );
  INVX2TS U1970 ( .A(n2012), .Y(n1668) );
  INVX2TS U1971 ( .A(\addr_calc/fir_read_calc/count[20] ), .Y(n1984) );
  INVX2TS U1972 ( .A(\addr_calc/fir_read_calc/count[9] ), .Y(n1899) );
  INVX2TS U1973 ( .A(\addr_calc/fir_read_calc/count[28] ), .Y(n1870) );
  BUFX3TS U1974 ( .A(\addr_calc/fir_read_calc/count[5] ), .Y(n1904) );
  INVX2TS U1975 ( .A(\addr_calc/fir_read_calc/count[29] ), .Y(n1841) );
  INVX2TS U1976 ( .A(\addr_calc/fir_read_calc/count[30] ), .Y(n1837) );
  INVX2TS U1977 ( .A(n2008), .Y(n1669) );
  INVX2TS U1978 ( .A(n2337), .Y(n2338) );
  INVX2TS U1979 ( .A(n2326), .Y(n2327) );
  INVX2TS U1980 ( .A(n2339), .Y(n2340) );
  INVX2TS U1981 ( .A(n2331), .Y(n2332) );
  CLKINVX1TS U1982 ( .A(n2314), .Y(n2315) );
  INVX1TS U1983 ( .A(n2486), .Y(n2488) );
  INVX1TS U1984 ( .A(n2415), .Y(n2418) );
  INVX1TS U1985 ( .A(n2439), .Y(n2441) );
  INVX1TS U1986 ( .A(n2447), .Y(n2450) );
  INVX1TS U1987 ( .A(n2467), .Y(n2469) );
  INVX1TS U1988 ( .A(n2490), .Y(n2493) );
  INVX1TS U1989 ( .A(n2497), .Y(n2500) );
  INVX1TS U1990 ( .A(n2419), .Y(n2422) );
  INVX1TS U1991 ( .A(n2451), .Y(n2454) );
  CLKINVX2TS U1992 ( .A(n2443), .Y(n2444) );
  INVX1TS U1993 ( .A(n2427), .Y(n2428) );
  INVX1TS U1994 ( .A(n2471), .Y(n1864) );
  INVX1TS U1995 ( .A(n2403), .Y(n2404) );
  INVX1TS U1996 ( .A(n2411), .Y(n2412) );
  INVX1TS U1997 ( .A(n2415), .Y(n2416) );
  INVX1TS U1998 ( .A(n2423), .Y(n2426) );
  INVX1TS U1999 ( .A(n2478), .Y(n2481) );
  INVX1TS U2000 ( .A(n2407), .Y(n2409) );
  INVX1TS U2001 ( .A(n2403), .Y(n2405) );
  INVX1TS U2002 ( .A(n2463), .Y(n2466) );
  INVX1TS U2003 ( .A(n2471), .Y(n2473) );
  INVX1TS U2004 ( .A(n2383), .Y(n2385) );
  INVX1TS U2005 ( .A(n2435), .Y(n2437) );
  INVX1TS U2006 ( .A(n2443), .Y(n2446) );
  INVX1TS U2007 ( .A(n2482), .Y(n2485) );
  INVX1TS U2008 ( .A(n2395), .Y(n2397) );
  INVX1TS U2009 ( .A(n2471), .Y(n2472) );
  INVX1TS U2010 ( .A(n2463), .Y(n2464) );
  INVX1TS U2011 ( .A(n2467), .Y(n2470) );
  INVX1TS U2012 ( .A(n2486), .Y(n2489) );
  CLKINVX2TS U2013 ( .A(n2486), .Y(n2487) );
  INVX1TS U2014 ( .A(n2375), .Y(n2378) );
  INVX2TS U2015 ( .A(n1757), .Y(n1760) );
  INVX2TS U2016 ( .A(n1758), .Y(n1763) );
  INVX3TS U2017 ( .A(n1757), .Y(n1761) );
  INVX3TS U2018 ( .A(n1704), .Y(n1749) );
  INVX3TS U2019 ( .A(n1745), .Y(n1671) );
  INVX2TS U2020 ( .A(n1704), .Y(n1748) );
  INVX4TS U2021 ( .A(n1701), .Y(n1753) );
  CLKINVX6TS U2022 ( .A(\addr_calc/fft_write_calc/counter/N38 ), .Y(n1675) );
  XNOR2X1TS U2023 ( .A(\add_x_19_0/n50 ), .B(\add_x_19_0/n4 ), .Y(
        \addr_calc/fft_read_addr[28] ) );
  XNOR2X1TS U2024 ( .A(\add_x_19_3/n50 ), .B(\add_x_19_3/n4 ), .Y(
        \addr_calc/fir_write_addr[28] ) );
  OR3X2TS U2025 ( .A(\data_cntl/N99 ), .B(n2808), .C(n2060), .Y(n1696) );
  INVX1TS U2026 ( .A(\add_x_19_3/n92 ), .Y(\add_x_19_3/n91 ) );
  AOI21X1TS U2027 ( .A0(\add_x_19_5/n69 ), .A1(\add_x_19_5/n61 ), .B0(
        \add_x_19_5/n62 ), .Y(\add_x_19_5/n60 ) );
  INVX1TS U2028 ( .A(\add_x_19_5/n134 ), .Y(\add_x_19_5/n133 ) );
  INVX1TS U2029 ( .A(\add_x_19_1/n134 ), .Y(\add_x_19_1/n133 ) );
  CLKINVX2TS U2030 ( .A(\add_x_19_2/n134 ), .Y(\add_x_19_2/n133 ) );
  INVX1TS U2031 ( .A(\add_x_19_3/n134 ), .Y(\add_x_19_3/n133 ) );
  CLKINVX2TS U2032 ( .A(\add_x_22_0/n42 ), .Y(\add_x_22_0/n41 ) );
  CLKINVX2TS U2033 ( .A(\add_x_22_1/n42 ), .Y(\add_x_22_1/n41 ) );
  CLKINVX2TS U2034 ( .A(\add_x_22_2/n42 ), .Y(\add_x_22_2/n41 ) );
  CLKINVX2TS U2035 ( .A(\add_x_22_3/n42 ), .Y(\add_x_22_3/n41 ) );
  CLKINVX2TS U2036 ( .A(\add_x_22_5/n42 ), .Y(\add_x_22_5/n41 ) );
  INVX2TS U2037 ( .A(\add_x_19_3/n113 ), .Y(n1676) );
  INVX1TS U2038 ( .A(\add_x_19_5/n72 ), .Y(\add_x_19_5/n70 ) );
  INVX1TS U2039 ( .A(\add_x_22_1/n59 ), .Y(\add_x_22_1/n58 ) );
  INVX1TS U2040 ( .A(\add_x_22_4/n59 ), .Y(\add_x_22_4/n58 ) );
  INVX1TS U2041 ( .A(\add_x_22_5/n59 ), .Y(\add_x_22_5/n58 ) );
  OAI21X1TS U2042 ( .A0(\addr_calc/fft_write_calc/counter/N43 ), .A1(n2796), 
        .B0(n2073), .Y(n2798) );
  INVX1TS U2043 ( .A(\add_x_22_3/n59 ), .Y(\add_x_22_3/n58 ) );
  INVX1TS U2044 ( .A(\add_x_22_0/n59 ), .Y(\add_x_22_0/n58 ) );
  AOI21X1TS U2045 ( .A0(\add_x_19_1/n73 ), .A1(\add_x_19_1/n46 ), .B0(
        \add_x_19_1/n47 ), .Y(\add_x_19_1/n45 ) );
  INVX1TS U2046 ( .A(\add_x_22_2/n59 ), .Y(\add_x_22_2/n58 ) );
  AOI21X1TS U2047 ( .A0(\add_x_19_3/n62 ), .A1(\add_x_19_3/n53 ), .B0(
        \add_x_19_3/n54 ), .Y(\add_x_19_3/n52 ) );
  INVX2TS U2048 ( .A(n936), .Y(n1830) );
  INVX1TS U2049 ( .A(\add_x_19_3/n73 ), .Y(\add_x_19_3/n71 ) );
  NAND2X2TS U2050 ( .A(n1787), .B(n2365), .Y(\DP_OP_159_297_3515/n1031 ) );
  CLKINVX2TS U2051 ( .A(\add_x_22_3/n94 ), .Y(\add_x_22_3/n93 ) );
  CLKINVX2TS U2052 ( .A(\add_x_22_4/n94 ), .Y(\add_x_22_4/n93 ) );
  CLKINVX2TS U2053 ( .A(\add_x_22_2/n94 ), .Y(\add_x_22_2/n93 ) );
  OAI21X1TS U2054 ( .A0(\add_x_19_3/n94 ), .A1(\add_x_19_3/n74 ), .B0(
        \add_x_19_3/n75 ), .Y(\add_x_19_3/n73 ) );
  CLKINVX2TS U2055 ( .A(\add_x_22_5/n94 ), .Y(\add_x_22_5/n93 ) );
  OAI21X1TS U2056 ( .A0(n2791), .A1(n2790), .B0(n2815), .Y(n2792) );
  CLKINVX2TS U2057 ( .A(\add_x_22_1/n94 ), .Y(\add_x_22_1/n93 ) );
  CLKINVX1TS U2058 ( .A(\add_x_19_0/n149 ), .Y(\add_x_19_0/n147 ) );
  CLKINVX1TS U2059 ( .A(\add_x_19_1/n149 ), .Y(\add_x_19_1/n147 ) );
  CLKINVX1TS U2060 ( .A(\add_x_19_2/n149 ), .Y(\add_x_19_2/n147 ) );
  CLKINVX1TS U2061 ( .A(\add_x_19_3/n149 ), .Y(\add_x_19_3/n147 ) );
  CLKINVX1TS U2062 ( .A(\add_x_19_5/n149 ), .Y(\add_x_19_5/n147 ) );
  INVX1TS U2063 ( .A(\add_x_19_5/n150 ), .Y(\add_x_19_5/n148 ) );
  INVX1TS U2064 ( .A(\add_x_19_4/n150 ), .Y(\add_x_19_4/n148 ) );
  CLKINVX1TS U2065 ( .A(\add_x_19_4/n149 ), .Y(\add_x_19_4/n147 ) );
  AOI21X1TS U2066 ( .A0(\add_x_19_4/n137 ), .A1(\add_x_19_4/n150 ), .B0(
        \add_x_19_4/n138 ), .Y(\add_x_19_4/n136 ) );
  INVX1TS U2067 ( .A(\add_x_22_5/n111 ), .Y(\add_x_22_5/n110 ) );
  INVX1TS U2068 ( .A(\add_x_22_3/n111 ), .Y(\add_x_22_3/n110 ) );
  AOI21X1TS U2069 ( .A0(\add_x_19_1/n95 ), .A1(\add_x_19_1/n104 ), .B0(
        \add_x_19_1/n96 ), .Y(\add_x_19_1/n94 ) );
  AOI21X1TS U2070 ( .A0(\add_x_19_3/n95 ), .A1(\add_x_19_3/n104 ), .B0(
        \add_x_19_3/n96 ), .Y(\add_x_19_3/n94 ) );
  INVX1TS U2071 ( .A(\add_x_19_1/n178 ), .Y(\add_x_19_1/n177 ) );
  AOI21X1TS U2072 ( .A0(\add_x_19_4/n76 ), .A1(\add_x_19_4/n85 ), .B0(
        \add_x_19_4/n77 ), .Y(\add_x_19_4/n75 ) );
  AOI21X1TS U2073 ( .A0(\add_x_19_0/n53 ), .A1(\add_x_19_0/n62 ), .B0(
        \add_x_19_0/n54 ), .Y(\add_x_19_0/n52 ) );
  INVX1TS U2074 ( .A(\add_x_22_0/n111 ), .Y(\add_x_22_0/n110 ) );
  INVX1TS U2075 ( .A(\add_x_22_4/n111 ), .Y(\add_x_22_4/n110 ) );
  CLKINVX1TS U2076 ( .A(\add_x_19_5/n151 ), .Y(\add_x_19_5/n214 ) );
  INVX1TS U2077 ( .A(\DP_OP_159_297_3515/n852 ), .Y(\DP_OP_159_297_3515/n928 )
         );
  OAI21X1TS U2078 ( .A0(\add_x_19_1/n151 ), .A1(\add_x_19_1/n155 ), .B0(
        \add_x_19_1/n152 ), .Y(\add_x_19_1/n150 ) );
  CLKINVX1TS U2079 ( .A(\add_x_19_0/n120 ), .Y(\add_x_19_0/n208 ) );
  CLKINVX1TS U2080 ( .A(\add_x_19_0/n97 ), .Y(\add_x_19_0/n204 ) );
  CLKINVX2TS U2081 ( .A(n2584), .Y(n2585) );
  CLKINVX1TS U2082 ( .A(\add_x_19_3/n97 ), .Y(\add_x_19_3/n204 ) );
  CLKINVX1TS U2083 ( .A(\add_x_19_4/n86 ), .Y(\add_x_19_4/n202 ) );
  OAI21X1TS U2084 ( .A0(\add_x_19_3/n105 ), .A1(\add_x_19_3/n111 ), .B0(
        \add_x_19_3/n106 ), .Y(\add_x_19_3/n104 ) );
  INVX1TS U2085 ( .A(\add_x_19_3/n120 ), .Y(\add_x_19_3/n208 ) );
  CLKINVX1TS U2086 ( .A(\add_x_19_1/n86 ), .Y(\add_x_19_1/n202 ) );
  CLKINVX1TS U2087 ( .A(\add_x_19_0/n86 ), .Y(\add_x_19_0/n202 ) );
  CLKINVX1TS U2088 ( .A(\add_x_19_0/n128 ), .Y(\add_x_19_0/n210 ) );
  CLKINVX1TS U2089 ( .A(\add_x_19_4/n105 ), .Y(\add_x_19_4/n206 ) );
  CLKINVX1TS U2090 ( .A(\add_x_19_5/n86 ), .Y(\add_x_19_5/n202 ) );
  INVX1TS U2091 ( .A(\add_x_19_4/n110 ), .Y(\add_x_19_4/n207 ) );
  INVX1TS U2092 ( .A(\add_x_19_4/n111 ), .Y(\add_x_19_4/n109 ) );
  INVX1TS U2093 ( .A(\add_x_22_0/n119 ), .Y(\add_x_22_0/n118 ) );
  CLKINVX1TS U2094 ( .A(\add_x_19_3/n86 ), .Y(\add_x_19_3/n202 ) );
  INVX1TS U2095 ( .A(\add_x_19_2/n110 ), .Y(\add_x_19_2/n207 ) );
  INVX1TS U2096 ( .A(\add_x_22_4/n119 ), .Y(\add_x_22_4/n118 ) );
  INVX1TS U2097 ( .A(\add_x_22_2/n111 ), .Y(\add_x_22_2/n110 ) );
  CLKINVX1TS U2098 ( .A(\add_x_19_1/n63 ), .Y(\add_x_19_1/n198 ) );
  INVX1TS U2099 ( .A(\add_x_22_1/n111 ), .Y(\add_x_22_1/n110 ) );
  CLKINVX1TS U2100 ( .A(\add_x_19_4/n66 ), .Y(\add_x_19_4/n199 ) );
  CLKINVX1TS U2101 ( .A(\add_x_19_3/n184 ), .Y(\add_x_19_3/n221 ) );
  CLKINVX1TS U2102 ( .A(\add_x_19_0/n63 ), .Y(\add_x_19_0/n198 ) );
  CLKINVX1TS U2103 ( .A(\add_x_19_5/n63 ), .Y(\add_x_19_5/n198 ) );
  INVX2TS U2104 ( .A(n2053), .Y(n2055) );
  INVX1TS U2105 ( .A(\add_x_19_4/n187 ), .Y(\add_x_19_4/n186 ) );
  INVX2TS U2106 ( .A(n2053), .Y(n2054) );
  NOR2X2TS U2107 ( .A(n1900), .B(n1980), .Y(\add_x_19_2/n151 ) );
  CLKAND2X2TS U2108 ( .A(n2342), .B(n2341), .Y(n2603) );
  CLKINVX1TS U2109 ( .A(\add_x_19_5/n181 ), .Y(\add_x_19_5/n220 ) );
  INVX1TS U2110 ( .A(\add_x_19_3/n175 ), .Y(\add_x_19_3/n219 ) );
  CLKINVX1TS U2111 ( .A(\add_x_19_3/n165 ), .Y(\add_x_19_3/n217 ) );
  INVX2TS U2112 ( .A(\add_x_22_1/n64 ), .Y(n1976) );
  INVX1TS U2113 ( .A(\add_x_22_2/n119 ), .Y(\add_x_22_2/n118 ) );
  INVX1TS U2114 ( .A(\add_x_22_3/n119 ), .Y(\add_x_22_3/n118 ) );
  CLKINVX1TS U2115 ( .A(\add_x_19_4/n139 ), .Y(\add_x_19_4/n212 ) );
  INVX1TS U2116 ( .A(\add_x_19_4/n144 ), .Y(\add_x_19_4/n213 ) );
  INVX1TS U2117 ( .A(\add_x_22_1/n119 ), .Y(\add_x_22_1/n118 ) );
  CLKINVX1TS U2118 ( .A(\add_x_19_1/n120 ), .Y(\add_x_19_1/n208 ) );
  CLKINVX1TS U2119 ( .A(\add_x_19_3/n154 ), .Y(\add_x_19_3/n215 ) );
  INVX2TS U2120 ( .A(\DP_OP_159_297_3515/n815 ), .Y(n2372) );
  NOR2X1TS U2121 ( .A(\add_x_19_1/n110 ), .B(\add_x_19_1/n105 ), .Y(
        \add_x_19_1/n103 ) );
  OAI21X1TS U2122 ( .A0(\add_x_19_1/n105 ), .A1(\add_x_19_1/n111 ), .B0(
        \add_x_19_1/n106 ), .Y(\add_x_19_1/n104 ) );
  NOR2X1TS U2123 ( .A(\add_x_19_2/n58 ), .B(\add_x_19_2/n55 ), .Y(
        \add_x_19_2/n53 ) );
  OAI21X1TS U2124 ( .A0(\add_x_19_4/n188 ), .A1(\add_x_19_4/n191 ), .B0(
        \add_x_19_4/n189 ), .Y(\add_x_19_4/n187 ) );
  INVX2TS U2125 ( .A(\DP_OP_159_297_3515/n877 ), .Y(n2362) );
  INVX1TS U2126 ( .A(\add_x_19_5/n144 ), .Y(\add_x_19_5/n213 ) );
  CLKINVX1TS U2127 ( .A(\add_x_19_4/n184 ), .Y(\add_x_19_4/n221 ) );
  INVX1TS U2128 ( .A(\add_x_19_3/n144 ), .Y(\add_x_19_3/n213 ) );
  CLKINVX1TS U2129 ( .A(\add_x_19_2/n139 ), .Y(\add_x_19_2/n212 ) );
  CLKINVX1TS U2130 ( .A(\DP_OP_159_297_3515/n943 ), .Y(
        \DP_OP_159_297_3515/n944 ) );
  CLKINVX1TS U2131 ( .A(\add_x_19_5/n128 ), .Y(\add_x_19_5/n210 ) );
  INVX2TS U2132 ( .A(n1562), .Y(n1678) );
  CLKINVX1TS U2133 ( .A(\add_x_19_1/n176 ), .Y(\add_x_19_1/n174 ) );
  CLKINVX1TS U2134 ( .A(\DP_OP_159_297_3515/n1026 ), .Y(
        \DP_OP_159_297_3515/n1025 ) );
  CLKINVX1TS U2135 ( .A(\add_x_19_3/n170 ), .Y(\add_x_19_3/n218 ) );
  CLKINVX1TS U2136 ( .A(\add_x_19_4/n165 ), .Y(\add_x_19_4/n217 ) );
  INVX2TS U2137 ( .A(\DP_OP_159_297_3515/n867 ), .Y(n2369) );
  CLKINVX1TS U2138 ( .A(\add_x_19_2/n154 ), .Y(\add_x_19_2/n215 ) );
  CLKINVX1TS U2139 ( .A(\add_x_19_0/n154 ), .Y(\add_x_19_0/n215 ) );
  CLKINVX1TS U2140 ( .A(\add_x_19_2/n128 ), .Y(\add_x_19_2/n210 ) );
  INVX1TS U2141 ( .A(\add_x_19_2/n175 ), .Y(\add_x_19_2/n219 ) );
  CLKINVX1TS U2142 ( .A(\add_x_19_2/n120 ), .Y(\add_x_19_2/n208 ) );
  INVX1TS U2143 ( .A(\add_x_19_3/n110 ), .Y(\add_x_19_3/n207 ) );
  INVX1TS U2144 ( .A(\add_x_19_0/n110 ), .Y(\add_x_19_0/n207 ) );
  INVX1TS U2145 ( .A(\add_x_19_3/n63 ), .Y(\add_x_19_3/n198 ) );
  CLKINVX1TS U2146 ( .A(\add_x_19_5/n105 ), .Y(\add_x_19_5/n206 ) );
  CLKINVX1TS U2147 ( .A(\add_x_19_2/n105 ), .Y(\add_x_19_2/n206 ) );
  INVX1TS U2148 ( .A(\add_x_19_5/n110 ), .Y(\add_x_19_5/n207 ) );
  CLKINVX2TS U2149 ( .A(\add_x_19_5/n111 ), .Y(\add_x_19_5/n109 ) );
  CLKINVX1TS U2150 ( .A(\add_x_19_1/n128 ), .Y(\add_x_19_1/n210 ) );
  CLKINVX1TS U2151 ( .A(\add_x_19_2/n97 ), .Y(\add_x_19_2/n204 ) );
  INVX1TS U2152 ( .A(\add_x_19_1/n110 ), .Y(\add_x_19_1/n207 ) );
  CLKINVX1TS U2153 ( .A(\add_x_19_4/n97 ), .Y(\add_x_19_4/n204 ) );
  INVX2TS U2154 ( .A(n2008), .Y(n2009) );
  INVX2TS U2155 ( .A(n1989), .Y(n1990) );
  INVX2TS U2156 ( .A(n2024), .Y(n2025) );
  INVX2TS U2157 ( .A(\add_x_22_2/n80 ), .Y(n1895) );
  INVX2TS U2158 ( .A(\add_x_22_2/n74 ), .Y(n1994) );
  CLKINVX1TS U2159 ( .A(n2070), .Y(n2072) );
  INVX2TS U2160 ( .A(\add_x_22_3/n71 ), .Y(n1880) );
  CLKINVX1TS U2161 ( .A(n2065), .Y(fir_enable) );
  INVX2TS U2162 ( .A(n2810), .Y(n2007) );
  INVX2TS U2163 ( .A(\add_x_22_3/n84 ), .Y(n1874) );
  INVX2TS U2164 ( .A(n1882), .Y(n1883) );
  INVX2TS U2165 ( .A(\add_x_22_3/n105 ), .Y(n1867) );
  INVX2TS U2166 ( .A(\add_x_22_3/n89 ), .Y(n1872) );
  INVX2TS U2167 ( .A(\add_x_22_3/n98 ), .Y(n1869) );
  INVX2TS U2168 ( .A(\add_x_22_3/n114 ), .Y(n1866) );
  INVX2TS U2169 ( .A(\add_x_22_4/n57 ), .Y(n1916) );
  INVX2TS U2170 ( .A(n2070), .Y(n2074) );
  INVX2TS U2171 ( .A(n1919), .Y(n1920) );
  INVX2TS U2172 ( .A(\add_x_22_5/n92 ), .Y(n2041) );
  INVX2TS U2173 ( .A(\add_x_22_2/n92 ), .Y(n1997) );
  INVX2TS U2174 ( .A(\add_x_22_2/n114 ), .Y(n1908) );
  INVX2TS U2175 ( .A(n1844), .Y(n1845) );
  INVX2TS U2176 ( .A(\add_x_22_5/n109 ), .Y(n1935) );
  INVX2TS U2177 ( .A(\add_x_22_5/n71 ), .Y(n1945) );
  INVX2TS U2178 ( .A(\add_x_22_5/n64 ), .Y(n1948) );
  INVX2TS U2179 ( .A(\add_x_22_5/n57 ), .Y(n1951) );
  INVX2TS U2180 ( .A(n1878), .Y(n1879) );
  INVX2TS U2181 ( .A(\add_x_22_5/n53 ), .Y(n1954) );
  INVX2TS U2182 ( .A(n1887), .Y(n1888) );
  INVX2TS U2183 ( .A(\add_x_22_2/n109 ), .Y(n1906) );
  INVX2TS U2184 ( .A(n2019), .Y(n2020) );
  INVX2TS U2185 ( .A(\add_x_22_2/n101 ), .Y(n2001) );
  INVX2TS U2186 ( .A(\add_x_22_5/n74 ), .Y(n2044) );
  INVX2TS U2187 ( .A(\add_x_22_5/n80 ), .Y(n1942) );
  INVX2TS U2188 ( .A(\add_x_22_3/n7 ), .Y(n1896) );
  INVX2TS U2189 ( .A(n1832), .Y(n1833) );
  INVX2TS U2190 ( .A(\add_x_22_5/n84 ), .Y(n1940) );
  INVX2TS U2191 ( .A(\add_x_22_2/n12 ), .Y(n1873) );
  INVX2TS U2192 ( .A(n1841), .Y(n1842) );
  INVX2TS U2193 ( .A(\add_x_22_2/n46 ), .Y(n1881) );
  INVX2TS U2194 ( .A(\add_x_22_2/n53 ), .Y(n1884) );
  INVX2TS U2195 ( .A(\add_x_22_2/n71 ), .Y(n1893) );
  INVX2TS U2196 ( .A(\add_x_22_5/n101 ), .Y(n2039) );
  INVX2TS U2197 ( .A(\add_x_22_2/n64 ), .Y(n1890) );
  INVX2TS U2198 ( .A(\add_x_22_1/n84 ), .Y(n1932) );
  INVX2TS U2199 ( .A(\addr_calc/fft_write_calc/count[15] ), .Y(
        \add_x_22_1/n64 ) );
  CLKINVX1TS U2200 ( .A(n2035), .Y(\addr_calc/fft_write_calc/counter/N43 ) );
  INVX2TS U2201 ( .A(\add_x_22_1/n71 ), .Y(n1927) );
  INVX1TS U2202 ( .A(\addr_calc/iir_read_calc/count[10] ), .Y(\add_x_22_4/n84 ) );
  CLKINVX1TS U2203 ( .A(\addr_calc/iir_read_calc/count[7] ), .Y(
        \add_x_22_4/n98 ) );
  INVX2TS U2204 ( .A(\add_x_22_1/n74 ), .Y(n2023) );
  INVX2TS U2205 ( .A(n1952), .Y(n1953) );
  INVX2TS U2206 ( .A(\add_x_22_0/n92 ), .Y(n2049) );
  INVX2TS U2207 ( .A(\add_x_22_0/n101 ), .Y(n2052) );
  INVX2TS U2208 ( .A(n2062), .Y(n2063) );
  CLKINVX1TS U2209 ( .A(\addr_calc/iir_read_calc/count[11] ), .Y(
        \add_x_22_4/n80 ) );
  INVX2TS U2210 ( .A(n1828), .Y(n1829) );
  CLKINVX1TS U2211 ( .A(n2022), .Y(\add_x_22_1/n67 ) );
  INVX2TS U2212 ( .A(n1852), .Y(n1853) );
  INVX1TS U2213 ( .A(n2552), .Y(\add_x_22_0/n109 ) );
  CLKINVX1TS U2214 ( .A(n1977), .Y(\add_x_22_0/n105 ) );
  CLKINVX4TS U2215 ( .A(n2057), .Y(n2058) );
  INVX2TS U2216 ( .A(n1855), .Y(n1856) );
  CLKINVX1TS U2217 ( .A(n1993), .Y(\add_x_22_3/n101 ) );
  INVX1TS U2218 ( .A(\addr_calc/fir_write_calc/count[4] ), .Y(
        \add_x_22_3/n109 ) );
  INVX1TS U2219 ( .A(n1943), .Y(n1944) );
  CLKINVX1TS U2220 ( .A(n1996), .Y(\add_x_22_3/n92 ) );
  INVX2TS U2221 ( .A(\add_x_22_4/n33 ), .Y(n2031) );
  INVX2TS U2222 ( .A(\add_x_22_1/n98 ), .Y(n1936) );
  INVX2TS U2223 ( .A(n1862), .Y(n1863) );
  INVX2TS U2224 ( .A(\add_x_22_1/n92 ), .Y(n2026) );
  INVX2TS U2225 ( .A(\add_x_22_1/n89 ), .Y(n1934) );
  INVX2TS U2226 ( .A(\add_x_22_4/n101 ), .Y(n2018) );
  INVX2TS U2227 ( .A(\add_x_22_1/n53 ), .Y(n1924) );
  CLKINVX1TS U2228 ( .A(\addr_calc/fir_read_calc/count[1] ), .Y(
        \add_x_22_2/n121 ) );
  INVX2TS U2229 ( .A(\add_x_22_0/n84 ), .Y(n1972) );
  CLKINVX1TS U2230 ( .A(\addr_calc/fir_read_calc/count[5] ), .Y(
        \add_x_22_2/n105 ) );
  INVX1TS U2231 ( .A(n1894), .Y(\add_x_22_3/n19 ) );
  INVX2TS U2232 ( .A(\add_x_22_0/n80 ), .Y(n1970) );
  CLKINVX1TS U2233 ( .A(n2065), .Y(n2069) );
  INVX2TS U2234 ( .A(n1968), .Y(n1969) );
  INVX2TS U2235 ( .A(n1839), .Y(n1840) );
  CLKINVX2TS U2236 ( .A(\add_x_22_4/n105 ), .Y(n2553) );
  INVX2TS U2237 ( .A(\add_x_22_3/n80 ), .Y(n1877) );
  INVX2TS U2238 ( .A(n1973), .Y(n1974) );
  CLKINVX1TS U2239 ( .A(\addr_calc/iir_write_calc/count[3] ), .Y(
        \add_x_22_5/n114 ) );
  NOR2X1TS U2240 ( .A(\addr_calc/iir_read_calc/count[28] ), .B(n2384), .Y(
        \add_x_19_4/n48 ) );
  NOR2X1TS U2241 ( .A(\addr_calc/iir_read_calc/count[19] ), .B(n2487), .Y(
        \add_x_19_4/n97 ) );
  NOR2X1TS U2242 ( .A(\addr_calc/iir_read_calc/count[26] ), .B(n2376), .Y(
        \add_x_19_4/n58 ) );
  NOR2X1TS U2243 ( .A(\addr_calc/fft_write_calc/count[23] ), .B(n2468), .Y(
        \add_x_19_1/n78 ) );
  NOR2X1TS U2244 ( .A(\addr_calc/fft_write_calc/count[26] ), .B(n2378), .Y(
        \add_x_19_1/n58 ) );
  NOR2X1TS U2245 ( .A(\addr_calc/fft_write_calc/count[28] ), .B(n2386), .Y(
        \add_x_19_1/n48 ) );
  NOR2X1TS U2246 ( .A(\addr_calc/fft_write_calc/count[16] ), .B(n2400), .Y(
        \add_x_19_1/n110 ) );
  NOR2X1TS U2247 ( .A(\addr_calc/fir_read_calc/count[4] ), .B(n2396), .Y(
        \add_x_19_2/n175 ) );
  NOR2X1TS U2248 ( .A(\addr_calc/iir_write_calc/count[22] ), .B(n2465), .Y(
        \add_x_19_5/n81 ) );
  NOR2X1TS U2249 ( .A(\addr_calc/iir_write_calc/count[26] ), .B(n2377), .Y(
        \add_x_19_5/n58 ) );
  INVX2TS U2250 ( .A(\DP_OP_159_297_3515/n950 ), .Y(n1679) );
  NOR2X1TS U2251 ( .A(\addr_calc/fir_write_calc/count[26] ), .B(n2376), .Y(
        \add_x_19_3/n58 ) );
  NOR2X1TS U2252 ( .A(\addr_calc/fft_read_calc/count[28] ), .B(n2385), .Y(
        \add_x_19_0/n48 ) );
  NOR2X1TS U2253 ( .A(\addr_calc/fir_write_calc/count[24] ), .B(n2462), .Y(
        \add_x_19_3/n66 ) );
  NOR2X1TS U2254 ( .A(\addr_calc/fft_read_calc/count[26] ), .B(n2376), .Y(
        \add_x_19_0/n58 ) );
  NOR2X1TS U2255 ( .A(\addr_calc/fir_write_calc/count[23] ), .B(n2468), .Y(
        \add_x_19_3/n78 ) );
  INVX2TS U2256 ( .A(n1456), .Y(n1680) );
  INVX2TS U2257 ( .A(\DP_OP_159_297_3515/n873 ), .Y(n1681) );
  OR2X1TS U2258 ( .A(\addr_calc/fir_write_calc/count[31] ), .B(n2381), .Y(
        n2630) );
  NOR2X1TS U2259 ( .A(\addr_calc/fir_write_calc/count[16] ), .B(n2401), .Y(
        \add_x_19_3/n110 ) );
  INVX2TS U2260 ( .A(\DP_OP_159_297_3515/n871 ), .Y(n1682) );
  BUFX3TS U2261 ( .A(\addr_calc/iir_read_calc/count[7] ), .Y(n1905) );
  INVX2TS U2262 ( .A(\addr_calc/fft_read_calc/count[9] ), .Y(\add_x_22_0/n89 )
         );
  CLKBUFX2TS U2263 ( .A(\addr_calc/fft_read_calc/count[4] ), .Y(n2552) );
  INVX2TS U2264 ( .A(\addr_calc/iir_write_calc/count[29] ), .Y(n1850) );
  INVX2TS U2265 ( .A(\addr_calc/fft_read_calc/count[8] ), .Y(\add_x_22_0/n92 )
         );
  INVX2TS U2266 ( .A(\addr_calc/fir_write_calc/count[23] ), .Y(
        \add_x_22_3/n30 ) );
  INVX2TS U2267 ( .A(\addr_calc/iir_write_calc/count[28] ), .Y(n1973) );
  INVX2TS U2268 ( .A(\addr_calc/fft_write_calc/count[12] ), .Y(
        \add_x_22_1/n74 ) );
  INVX2TS U2269 ( .A(n1843), .Y(n1684) );
  INVX2TS U2270 ( .A(n1907), .Y(n1685) );
  INVX2TS U2271 ( .A(\addr_calc/fir_write_calc/count[26] ), .Y(
        \add_x_22_3/n15 ) );
  INVX2TS U2272 ( .A(\addr_calc/fft_read_calc/count[18] ), .Y(\add_x_22_0/n49 ) );
  INVX2TS U2273 ( .A(\addr_calc/iir_read_calc/count[28] ), .Y(\add_x_22_4/n7 )
         );
  INVX2TS U2274 ( .A(\addr_calc/fft_write_calc/count[13] ), .Y(
        \add_x_22_1/n71 ) );
  INVX2TS U2275 ( .A(\addr_calc/iir_read_calc/count[29] ), .Y(n1839) );
  INVX2TS U2276 ( .A(\addr_calc/iir_write_calc/count[23] ), .Y(n1964) );
  INVX2TS U2277 ( .A(\addr_calc/fft_read_calc/count[10] ), .Y(\add_x_22_0/n84 ) );
  INVX2TS U2278 ( .A(n1923), .Y(n1687) );
  INVX2TS U2279 ( .A(\addr_calc/fft_read_calc/count[11] ), .Y(\add_x_22_0/n80 ) );
  INVX2TS U2280 ( .A(\addr_calc/fft_write_calc/count[17] ), .Y(
        \add_x_22_1/n53 ) );
  INVX2TS U2281 ( .A(\addr_calc/iir_write_calc/count[19] ), .Y(n1957) );
  INVX2TS U2282 ( .A(\addr_calc/iir_write_calc/count[24] ), .Y(n2050) );
  INVX2TS U2283 ( .A(\addr_calc/iir_read_calc/count[17] ), .Y(n1919) );
  INVX2TS U2284 ( .A(\addr_calc/fir_write_calc/count[11] ), .Y(
        \add_x_22_3/n80 ) );
  INVX2TS U2285 ( .A(\addr_calc/fir_write_calc/count[5] ), .Y(
        \add_x_22_3/n105 ) );
  INVX2TS U2286 ( .A(n1971), .Y(n1688) );
  INVX2TS U2287 ( .A(\addr_calc/iir_read_calc/count[23] ), .Y(\add_x_22_4/n30 ) );
  INVX2TS U2288 ( .A(\addr_calc/fft_read_calc/count[31] ), .Y(n1855) );
  INVX2TS U2289 ( .A(\addr_calc/iir_read_calc/count[13] ), .Y(\add_x_22_4/n71 ) );
  INVX2TS U2290 ( .A(n2814), .Y(n2065) );
  INVX2TS U2291 ( .A(n2815), .Y(n2062) );
  INVX2TS U2292 ( .A(\addr_calc/iir_read_calc/count[0] ), .Y(n2786) );
  INVX2TS U2293 ( .A(\addr_calc/iir_write_calc/count[0] ), .Y(n2791) );
  INVX2TS U2294 ( .A(\addr_calc/iir_read_calc/count[8] ), .Y(\add_x_22_4/n92 )
         );
  INVX2TS U2295 ( .A(\addr_calc/fft_write_calc/count[23] ), .Y(
        \add_x_22_1/n30 ) );
  INVX2TS U2296 ( .A(\addr_calc/fft_read_calc/count[22] ), .Y(n2040) );
  INVX2TS U2297 ( .A(\addr_calc/fft_write_calc/count[3] ), .Y(
        \add_x_22_1/n114 ) );
  INVX2TS U2298 ( .A(\addr_calc/fft_read_calc/count[27] ), .Y(n1943) );
  INVX2TS U2299 ( .A(\addr_calc/fft_read_calc/count[28] ), .Y(\add_x_22_0/n7 )
         );
  INVX2TS U2300 ( .A(\addr_calc/fft_write_calc/count[7] ), .Y(\add_x_22_1/n98 ) );
  INVX2TS U2301 ( .A(\addr_calc/fft_read_calc/count[29] ), .Y(n1862) );
  INVX2TS U2302 ( .A(\addr_calc/fft_write_calc/count[8] ), .Y(\add_x_22_1/n92 ) );
  INVX2TS U2303 ( .A(\addr_calc/fft_write_calc/count[9] ), .Y(\add_x_22_1/n89 ) );
  INVX2TS U2304 ( .A(\addr_calc/fft_write_calc/count[10] ), .Y(
        \add_x_22_1/n84 ) );
  INVX2TS U2305 ( .A(\addr_calc/fft_write_calc/count[26] ), .Y(
        \add_x_22_1/n15 ) );
  INVX2TS U2306 ( .A(\addr_calc/fir_read_calc/count[17] ), .Y(\add_x_22_2/n53 ) );
  INVX2TS U2307 ( .A(\addr_calc/fir_read_calc/count[3] ), .Y(\add_x_22_2/n114 ) );
  INVX2TS U2308 ( .A(\addr_calc/fir_read_calc/count[8] ), .Y(\add_x_22_2/n92 )
         );
  INVX2TS U2309 ( .A(\addr_calc/iir_write_calc/count[15] ), .Y(
        \add_x_22_5/n64 ) );
  INVX2TS U2310 ( .A(\addr_calc/fir_read_calc/count[4] ), .Y(\add_x_22_2/n109 ) );
  INVX2TS U2311 ( .A(\addr_calc/iir_write_calc/count[9] ), .Y(\add_x_22_5/n89 ) );
  INVX2TS U2312 ( .A(\addr_calc/iir_write_calc/count[26] ), .Y(
        \add_x_22_5/n15 ) );
  INVX2TS U2313 ( .A(\addr_calc/iir_write_calc/count[11] ), .Y(
        \add_x_22_5/n80 ) );
  INVX2TS U2314 ( .A(\addr_calc/fir_read_calc/count[19] ), .Y(\add_x_22_2/n46 ) );
  INVX2TS U2315 ( .A(\addr_calc/fir_read_calc/count[15] ), .Y(\add_x_22_2/n64 ) );
  INVX2TS U2316 ( .A(\addr_calc/iir_write_calc/count[8] ), .Y(\add_x_22_5/n92 ) );
  INVX2TS U2317 ( .A(\addr_calc/fir_read_calc/count[12] ), .Y(\add_x_22_2/n74 ) );
  INVX2TS U2318 ( .A(\addr_calc/fir_read_calc/count[11] ), .Y(\add_x_22_2/n80 ) );
  INVX2TS U2319 ( .A(\addr_calc/fir_write_calc/count[7] ), .Y(\add_x_22_3/n98 ) );
  INVX2TS U2320 ( .A(\addr_calc/fft_write_calc/count[31] ), .Y(n1844) );
  INVX2TS U2321 ( .A(\addr_calc/fir_write_calc/count[9] ), .Y(\add_x_22_3/n89 ) );
  INVX2TS U2322 ( .A(n1981), .Y(n1691) );
  INVX2TS U2323 ( .A(\addr_calc/fft_write_calc/count[28] ), .Y(\add_x_22_1/n7 ) );
  INVX2TS U2324 ( .A(\addr_calc/iir_write_calc/count[16] ), .Y(
        \add_x_22_5/n57 ) );
  INVX2TS U2325 ( .A(\addr_calc/fft_write_calc/count[11] ), .Y(n1930) );
  INVX2TS U2326 ( .A(\addr_calc/fft_write_calc/count[29] ), .Y(n1852) );
  INVX2TS U2327 ( .A(\addr_calc/fir_read_calc/count[24] ), .Y(n1982) );
  INVX2TS U2328 ( .A(\addr_calc/fir_write_calc/count[29] ), .Y(n1832) );
  INVX2TS U2329 ( .A(\addr_calc/iir_write_calc/count[10] ), .Y(
        \add_x_22_5/n84 ) );
  INVX2TS U2330 ( .A(\addr_calc/fir_write_calc/count[27] ), .Y(n1834) );
  INVX2TS U2331 ( .A(\addr_calc/iir_write_calc/count[1] ), .Y(
        \add_x_22_5/n121 ) );
  INVX2TS U2332 ( .A(\addr_calc/fir_write_calc/count[28] ), .Y(\add_x_22_3/n7 ) );
  INVX2TS U2333 ( .A(\addr_calc/fir_write_calc/count[13] ), .Y(
        \add_x_22_3/n71 ) );
  INVX2TS U2334 ( .A(\addr_calc/fir_read_calc/count[13] ), .Y(\add_x_22_2/n71 ) );
  INVX1TS U2335 ( .A(n2151), .Y(n2152) );
  INVX1TS U2336 ( .A(n2159), .Y(n2160) );
  CLKINVX2TS U2337 ( .A(n2335), .Y(n2336) );
  CLKINVX2TS U2338 ( .A(n2503), .Y(n2504) );
  CLKINVX2TS U2339 ( .A(n2501), .Y(n2502) );
  CLKINVX2TS U2340 ( .A(n2505), .Y(n2506) );
  INVX1TS U2341 ( .A(n2291), .Y(n2292) );
  INVX1TS U2342 ( .A(n2201), .Y(n2202) );
  INVX1TS U2343 ( .A(n2279), .Y(n2280) );
  CLKINVX2TS U2344 ( .A(n2351), .Y(n2352) );
  INVX1TS U2345 ( .A(n2241), .Y(n2242) );
  INVX1TS U2346 ( .A(n2455), .Y(n2457) );
  INVX1TS U2347 ( .A(n2247), .Y(n2248) );
  CLKINVX2TS U2348 ( .A(n2309), .Y(n2310) );
  CLKINVX2TS U2349 ( .A(n2355), .Y(n2356) );
  CLKINVX1TS U2350 ( .A(n1798), .Y(n1799) );
  INVX1TS U2351 ( .A(n2163), .Y(n2164) );
  CLKINVX2TS U2352 ( .A(n2517), .Y(n2518) );
  CLKINVX1TS U2353 ( .A(n1804), .Y(n1805) );
  CLKINVX2TS U2354 ( .A(n2519), .Y(n2520) );
  INVX1TS U2355 ( .A(n2243), .Y(n2244) );
  CLKINVX2TS U2356 ( .A(n2533), .Y(n2534) );
  INVX1TS U2357 ( .A(n2197), .Y(n2198) );
  CLKINVX1TS U2358 ( .A(n1800), .Y(n1801) );
  INVX1TS U2359 ( .A(n2205), .Y(n2206) );
  INVX1TS U2360 ( .A(n2287), .Y(n2288) );
  INVX1TS U2361 ( .A(n2283), .Y(n2284) );
  CLKINVX2TS U2362 ( .A(n2535), .Y(n2536) );
  INVX1TS U2363 ( .A(n2155), .Y(n2156) );
  INVX1TS U2364 ( .A(n2119), .Y(n2120) );
  INVX1TS U2365 ( .A(n2115), .Y(n2116) );
  CLKINVX2TS U2366 ( .A(n2539), .Y(n2540) );
  INVX1TS U2367 ( .A(n2399), .Y(n2402) );
  INVX1TS U2368 ( .A(n2271), .Y(n2272) );
  INVX1TS U2369 ( .A(n2233), .Y(n2234) );
  INVX1TS U2370 ( .A(n2127), .Y(n2128) );
  INVX1TS U2371 ( .A(n2431), .Y(n2432) );
  CLKINVX2TS U2372 ( .A(n2345), .Y(n2346) );
  INVX1TS U2373 ( .A(n2143), .Y(n2144) );
  INVX1TS U2374 ( .A(n2217), .Y(n2218) );
  CLKINVX2TS U2375 ( .A(n2509), .Y(n2510) );
  INVX1TS U2376 ( .A(n2267), .Y(n2268) );
  CLKINVX2TS U2377 ( .A(n2525), .Y(n2526) );
  INVX1TS U2378 ( .A(n2139), .Y(n2140) );
  INVX1TS U2379 ( .A(n2415), .Y(n2417) );
  INVX1TS U2380 ( .A(n2255), .Y(n2256) );
  CLKINVX2TS U2381 ( .A(n2541), .Y(n2542) );
  INVX1TS U2382 ( .A(n2407), .Y(n2408) );
  INVX1TS U2383 ( .A(n2221), .Y(n2222) );
  CLKINVX2TS U2384 ( .A(n2547), .Y(n2548) );
  CLKINVX2TS U2385 ( .A(n2349), .Y(n2350) );
  INVX1TS U2386 ( .A(n2263), .Y(n2264) );
  CLKINVX2TS U2387 ( .A(n2531), .Y(n2532) );
  INVX1TS U2388 ( .A(n2229), .Y(n2230) );
  CLKINVX2TS U2389 ( .A(n2515), .Y(n2516) );
  INVX1TS U2390 ( .A(n2135), .Y(n2136) );
  INVX1TS U2391 ( .A(n1816), .Y(n1817) );
  CLKINVX2TS U2392 ( .A(n2357), .Y(n2358) );
  CLKINVX2TS U2393 ( .A(n2511), .Y(n2512) );
  INVX1TS U2394 ( .A(n2423), .Y(n2425) );
  CLKINVX2TS U2395 ( .A(n2545), .Y(n2546) );
  INVX1TS U2396 ( .A(n2131), .Y(n2132) );
  INVX1TS U2397 ( .A(n2225), .Y(n2226) );
  CLKINVX2TS U2398 ( .A(n2529), .Y(n2530) );
  CLKINVX2TS U2399 ( .A(n2527), .Y(n2528) );
  INVX1TS U2400 ( .A(n1808), .Y(n1809) );
  CLKINVX2TS U2401 ( .A(n2513), .Y(n2514) );
  CLKINVX2TS U2402 ( .A(n2353), .Y(n2354) );
  INVX1TS U2403 ( .A(n2259), .Y(n2260) );
  INVX1TS U2404 ( .A(n2209), .Y(n2210) );
  CLKINVX2TS U2405 ( .A(n2521), .Y(n2522) );
  INVX1TS U2406 ( .A(n2237), .Y(n2238) );
  CLKINVX2TS U2407 ( .A(n2537), .Y(n2538) );
  INVX1TS U2408 ( .A(n2275), .Y(n2276) );
  INVX1TS U2409 ( .A(n2123), .Y(n2124) );
  CLKINVX2TS U2410 ( .A(n2347), .Y(n2348) );
  INVX1TS U2411 ( .A(n2147), .Y(n2148) );
  CLKINVX2TS U2412 ( .A(n2507), .Y(n2508) );
  INVX1TS U2413 ( .A(n2431), .Y(n2433) );
  INVX1TS U2414 ( .A(n2387), .Y(n2390) );
  INVX1TS U2415 ( .A(n2251), .Y(n2252) );
  CLKINVX2TS U2416 ( .A(n2523), .Y(n2524) );
  INVX1TS U2417 ( .A(n2213), .Y(n2214) );
  INVX1TS U2418 ( .A(n2478), .Y(n2479) );
  INVX1TS U2419 ( .A(n2497), .Y(n2499) );
  CLKINVX2TS U2420 ( .A(n2543), .Y(n2544) );
  INVX1TS U2421 ( .A(n2223), .Y(n2224) );
  INVX1TS U2422 ( .A(n2285), .Y(n2286) );
  INVX1TS U2423 ( .A(n2474), .Y(n2477) );
  INVX1TS U2424 ( .A(n2399), .Y(n2400) );
  INVX1TS U2425 ( .A(n2261), .Y(n2262) );
  INVX2TS U2426 ( .A(n2328), .Y(n2329) );
  INVX1TS U2427 ( .A(n2199), .Y(n2200) );
  INVX1TS U2428 ( .A(n2474), .Y(n2476) );
  INVX1TS U2429 ( .A(n2399), .Y(n2401) );
  INVX1TS U2430 ( .A(n2161), .Y(n2162) );
  INVX1TS U2431 ( .A(n2435), .Y(n2436) );
  INVX1TS U2432 ( .A(n2133), .Y(n2134) );
  INVX1TS U2433 ( .A(n2478), .Y(n2480) );
  INVX1TS U2434 ( .A(n2077), .Y(n2078) );
  INVX1TS U2435 ( .A(n2289), .Y(n2290) );
  INVX1TS U2436 ( .A(n2098), .Y(n2099) );
  INVX1TS U2437 ( .A(n2431), .Y(n2434) );
  INVX1TS U2438 ( .A(n2227), .Y(n2228) );
  INVX1TS U2439 ( .A(n2195), .Y(n2196) );
  INVX1TS U2440 ( .A(n2179), .Y(n2180) );
  INVX1TS U2441 ( .A(n2109), .Y(n2110) );
  INVX1TS U2442 ( .A(n2379), .Y(n2380) );
  INVX1TS U2443 ( .A(n2165), .Y(n2166) );
  INVX1TS U2444 ( .A(n2391), .Y(n2392) );
  INVX2TS U2445 ( .A(n2322), .Y(n2323) );
  INVX1TS U2446 ( .A(n2111), .Y(n2112) );
  INVX1TS U2447 ( .A(n2447), .Y(n2448) );
  INVX1TS U2448 ( .A(n2257), .Y(n2258) );
  INVX1TS U2449 ( .A(n2451), .Y(n2453) );
  INVX1TS U2450 ( .A(n2439), .Y(n2442) );
  INVX1TS U2451 ( .A(n2293), .Y(n2294) );
  INVX1TS U2452 ( .A(n2395), .Y(n2396) );
  INVX1TS U2453 ( .A(n2447), .Y(n2449) );
  INVX1TS U2454 ( .A(n2129), .Y(n2130) );
  INVX1TS U2455 ( .A(n2482), .Y(n2483) );
  INVX1TS U2456 ( .A(n2083), .Y(n2084) );
  INVX1TS U2457 ( .A(n2273), .Y(n2274) );
  INVX1TS U2458 ( .A(n2211), .Y(n2212) );
  INVX1TS U2459 ( .A(n2145), .Y(n2146) );
  INVX1TS U2460 ( .A(n2102), .Y(n2103) );
  INVX1TS U2461 ( .A(n2149), .Y(n2150) );
  INVX1TS U2462 ( .A(n2395), .Y(n2398) );
  INVX1TS U2463 ( .A(n2075), .Y(n2076) );
  INVX1TS U2464 ( .A(n2215), .Y(n2216) );
  INVX1TS U2465 ( .A(n2277), .Y(n2278) );
  INVX2TS U2466 ( .A(n2333), .Y(n2334) );
  INVX1TS U2467 ( .A(n2269), .Y(n2270) );
  INVX1TS U2468 ( .A(n2089), .Y(n2090) );
  INVX2TS U2469 ( .A(n2316), .Y(n2317) );
  INVX1TS U2470 ( .A(n2427), .Y(n2430) );
  INVX1TS U2471 ( .A(n2207), .Y(n2208) );
  INVX1TS U2472 ( .A(n2141), .Y(n2142) );
  INVX1TS U2473 ( .A(n2153), .Y(n2154) );
  CLKINVX1TS U2474 ( .A(n2320), .Y(n2321) );
  CLKINVX1TS U2475 ( .A(n2318), .Y(n2319) );
  INVX1TS U2476 ( .A(n2403), .Y(n2406) );
  INVX1TS U2477 ( .A(n2219), .Y(n2220) );
  INVX1TS U2478 ( .A(n2281), .Y(n2282) );
  INVX1TS U2479 ( .A(n2091), .Y(n2092) );
  INVX1TS U2480 ( .A(n2203), .Y(n2204) );
  INVX1TS U2481 ( .A(n2137), .Y(n2138) );
  INVX1TS U2482 ( .A(n2157), .Y(n2158) );
  INVX1TS U2483 ( .A(n2307), .Y(n2308) );
  INVX1TS U2484 ( .A(n2474), .Y(n2475) );
  INVX1TS U2485 ( .A(n2235), .Y(n2236) );
  INVX1TS U2486 ( .A(n2303), .Y(n2304) );
  INVX1TS U2487 ( .A(n2079), .Y(n2080) );
  INVX1TS U2488 ( .A(n2301), .Y(n2302) );
  CLKINVX2TS U2489 ( .A(n2497), .Y(n2498) );
  INVX1TS U2490 ( .A(n2175), .Y(n2176) );
  INVX1TS U2491 ( .A(n2411), .Y(n2413) );
  INVX1TS U2492 ( .A(n2249), .Y(n2250) );
  INVX1TS U2493 ( .A(n2185), .Y(n2186) );
  INVX1TS U2494 ( .A(n2383), .Y(n2384) );
  INVX1TS U2495 ( .A(n2183), .Y(n2184) );
  INVX1TS U2496 ( .A(n2379), .Y(n2382) );
  INVX1TS U2497 ( .A(n2085), .Y(n2086) );
  INVX1TS U2498 ( .A(n2387), .Y(n2389) );
  INVX1TS U2499 ( .A(n2121), .Y(n2122) );
  INVX1TS U2500 ( .A(n2299), .Y(n2300) );
  INVX1TS U2501 ( .A(n2094), .Y(n2095) );
  INVX1TS U2502 ( .A(n2387), .Y(n2388) );
  INVX1TS U2503 ( .A(n1802), .Y(n1803) );
  INVX1TS U2504 ( .A(n2177), .Y(n2178) );
  INVX1TS U2505 ( .A(n2459), .Y(n2461) );
  INVX1TS U2506 ( .A(n2455), .Y(n2456) );
  INVX2TS U2507 ( .A(n2324), .Y(n2325) );
  INVX1TS U2508 ( .A(n2171), .Y(n2172) );
  INVX1TS U2509 ( .A(n2239), .Y(n2240) );
  INVX1TS U2510 ( .A(n2305), .Y(n2306) );
  INVX1TS U2511 ( .A(n2455), .Y(n2458) );
  INVX1TS U2512 ( .A(n2189), .Y(n2190) );
  INVX1TS U2513 ( .A(n2113), .Y(n2114) );
  INVX1TS U2514 ( .A(n2245), .Y(n2246) );
  INVX1TS U2515 ( .A(n2295), .Y(n2296) );
  INVX1TS U2516 ( .A(n2167), .Y(n2168) );
  INVX1TS U2517 ( .A(n2383), .Y(n2386) );
  CLKINVX2TS U2518 ( .A(n2359), .Y(n2360) );
  INVX1TS U2519 ( .A(n2193), .Y(n2194) );
  INVX1TS U2520 ( .A(n2117), .Y(n2118) );
  INVX1TS U2521 ( .A(n2265), .Y(n2266) );
  INVX1TS U2522 ( .A(n2104), .Y(n2105) );
  INVX1TS U2523 ( .A(n2081), .Y(n2082) );
  INVX1TS U2524 ( .A(n2100), .Y(n2101) );
  INVX1TS U2525 ( .A(n2459), .Y(n2460) );
  INVX1TS U2526 ( .A(n2375), .Y(n2376) );
  INVX1TS U2527 ( .A(n2169), .Y(n2170) );
  INVX1TS U2528 ( .A(n2096), .Y(n2097) );
  INVX1TS U2529 ( .A(n2106), .Y(n2107) );
  INVX1TS U2530 ( .A(n2297), .Y(n2298) );
  INVX1TS U2531 ( .A(n2253), .Y(n2254) );
  INVX1TS U2532 ( .A(n2459), .Y(n2462) );
  INVX1TS U2533 ( .A(n2443), .Y(n2445) );
  INVX1TS U2534 ( .A(n2231), .Y(n2232) );
  INVX1TS U2535 ( .A(n2187), .Y(n2188) );
  INVX1TS U2536 ( .A(n2467), .Y(n2468) );
  INVX1TS U2537 ( .A(n2490), .Y(n2491) );
  INVX1TS U2538 ( .A(n2379), .Y(n2381) );
  INVX1TS U2539 ( .A(n2087), .Y(n2088) );
  INVX1TS U2540 ( .A(n2181), .Y(n2182) );
  INVX1TS U2541 ( .A(n2463), .Y(n2465) );
  INVX1TS U2542 ( .A(n2173), .Y(n2174) );
  INVX1TS U2543 ( .A(n2191), .Y(n2192) );
  INVX1TS U2544 ( .A(n2125), .Y(n2126) );
  INVX2TS U2545 ( .A(n2407), .Y(n2410) );
  INVX2TS U2546 ( .A(n2423), .Y(n2424) );
  XOR2X4TS U2547 ( .A(\DP_OP_159_297_3515/n989 ), .B(n2361), .Y(n2615) );
  AO22X4TS U2548 ( .A0(n1761), .A1(\addr_calc/fir_write_calc/counter/N57 ), 
        .B0(n1269), .B1(\addr_calc/fir_write_calc/count[14] ), .Y(n1116) );
  INVX2TS U2549 ( .A(n1946), .Y(n1947) );
  NOR2X2TS U2550 ( .A(\DP_OP_158_296_6262/n322 ), .B(\DP_OP_158_296_6262/n329 ), .Y(\DP_OP_158_296_6262/n320 ) );
  BUFX4TS U2551 ( .A(n2661), .Y(n2659) );
  XOR2X4TS U2552 ( .A(n1736), .B(n1678), .Y(n2602) );
  NOR2BX4TS U2553 ( .AN(n1692), .B(\DP_OP_159_297_3515/n650 ), .Y(
        \DP_OP_159_297_3515/n648 ) );
  XOR2X4TS U2554 ( .A(n2616), .B(n1948), .Y(n1692) );
  OAI21X2TS U2555 ( .A0(\add_x_19_4/n60 ), .A1(\add_x_19_4/n58 ), .B0(
        \add_x_19_4/n59 ), .Y(\add_x_19_4/n57 ) );
  AOI21X4TS U2556 ( .A0(\add_x_19_4/n69 ), .A1(\add_x_19_4/n61 ), .B0(
        \add_x_19_4/n62 ), .Y(\add_x_19_4/n60 ) );
  NOR2X4TS U2557 ( .A(\DP_OP_159_297_3515/n625 ), .B(\DP_OP_159_297_3515/n638 ), .Y(\DP_OP_159_297_3515/n623 ) );
  NOR2X4TS U2558 ( .A(\DP_OP_159_297_3515/n589 ), .B(\DP_OP_159_297_3515/n646 ), .Y(\DP_OP_159_297_3515/n587 ) );
  NAND2X4TS U2559 ( .A(\DP_OP_159_297_3515/n591 ), .B(
        \DP_OP_159_297_3515/n623 ), .Y(\DP_OP_159_297_3515/n589 ) );
  XNOR2X2TS U2560 ( .A(n2622), .B(n2041), .Y(\DP_OP_159_297_3515/n730 ) );
  AO22X4TS U2561 ( .A0(n1762), .A1(\addr_calc/fir_write_calc/counter/N65 ), 
        .B0(n1268), .B1(\addr_calc/fir_write_calc/count[22] ), .Y(n1108) );
  NOR2X2TS U2562 ( .A(\addr_calc/fir_write_calc/count[25] ), .B(n2493), .Y(
        \add_x_19_3/n63 ) );
  NOR2X2TS U2563 ( .A(\DP_OP_158_296_6262/n148 ), .B(\DP_OP_158_296_6262/n133 ), .Y(\DP_OP_158_296_6262/n131 ) );
  INVX2TS U2564 ( .A(n1719), .Y(n1724) );
  NOR2X4TS U2565 ( .A(\DP_OP_159_297_3515/n726 ), .B(\DP_OP_159_297_3515/n690 ), .Y(\DP_OP_159_297_3515/n688 ) );
  AND2X8TS U2566 ( .A(\DP_OP_159_297_3515/n587 ), .B(\DP_OP_159_297_3515/n688 ), .Y(n1780) );
  NAND2X2TS U2567 ( .A(n1791), .B(\DP_OP_159_297_3515/n914 ), .Y(
        \DP_OP_159_297_3515/n913 ) );
  NOR2X1TS U2568 ( .A(\DP_OP_158_296_6262/n1863 ), .B(n1664), .Y(
        \DP_OP_158_296_6262/n1855 ) );
  AO22X4TS U2569 ( .A0(n1760), .A1(\addr_calc/fir_write_calc/counter/N45 ), 
        .B0(n1270), .B1(n1990), .Y(n1128) );
  INVX2TS U2570 ( .A(n1758), .Y(n1764) );
  NAND2X2TS U2571 ( .A(n1792), .B(\DP_OP_159_297_3515/n935 ), .Y(
        \DP_OP_159_297_3515/n934 ) );
  XNOR2X4TS U2572 ( .A(\add_x_19_4/n99 ), .B(\add_x_19_4/n13 ), .Y(
        \addr_calc/iir_read_addr[19] ) );
  INVX2TS U2573 ( .A(\addr_calc/iir_write_calc/count[13] ), .Y(
        \add_x_22_5/n71 ) );
  XOR2X4TS U2574 ( .A(n1698), .B(\DP_OP_158_296_6262/n1897 ), .Y(n1697) );
  NOR4X1TS U2575 ( .A(n2076), .B(n2090), .C(n907), .D(n908), .Y(n906) );
  XOR2X4TS U2576 ( .A(\DP_OP_159_297_3515/n955 ), .B(n1679), .Y(n1699) );
  AO22X4TS U2577 ( .A0(n1822), .A1(\addr_calc/fir_read_calc/counter/N52 ), 
        .B0(n1672), .B1(\addr_calc/fir_read_calc/count[9] ), .Y(n1089) );
  AO22X4TS U2578 ( .A0(n1827), .A1(\addr_calc/fir_read_calc/counter/N63 ), 
        .B0(n1672), .B1(\addr_calc/fir_read_calc/count[20] ), .Y(n1078) );
  NOR2X4TS U2579 ( .A(\DP_OP_159_297_3515/n685 ), .B(\DP_OP_159_297_3515/n674 ), .Y(\DP_OP_159_297_3515/n672 ) );
  AO22X4TS U2580 ( .A0(n1755), .A1(\addr_calc/fft_read_calc/counter/N71 ), 
        .B0(n2659), .B1(n2559), .Y(n1006) );
  AO22X4TS U2581 ( .A0(n1749), .A1(\addr_calc/fft_read_calc/counter/N50 ), 
        .B0(n2655), .B1(n1666), .Y(n1027) );
  XNOR2X4TS U2582 ( .A(n2618), .B(n1945), .Y(\DP_OP_159_297_3515/n685 ) );
  AO22X4TS U2583 ( .A0(n1753), .A1(\addr_calc/fft_read_calc/counter/N63 ), 
        .B0(n1475), .B1(n2572), .Y(n1014) );
  CLKINVX3TS U2584 ( .A(n1782), .Y(n1792) );
  AO22X4TS U2585 ( .A0(n1750), .A1(\addr_calc/fft_read_calc/counter/N56 ), 
        .B0(n2657), .B1(\addr_calc/fft_read_calc/count[13] ), .Y(n1021) );
  AO22X4TS U2586 ( .A0(n1755), .A1(\addr_calc/fft_read_calc/counter/N57 ), 
        .B0(n2657), .B1(\addr_calc/fft_read_calc/count[14] ), .Y(n1020) );
  BUFX3TS U2587 ( .A(n2660), .Y(n2658) );
  AO22X4TS U2588 ( .A0(n1753), .A1(\addr_calc/fft_read_calc/counter/N55 ), 
        .B0(n2657), .B1(\addr_calc/fft_read_calc/count[12] ), .Y(n1022) );
  AO22X4TS U2589 ( .A0(n1750), .A1(\addr_calc/fft_read_calc/counter/N65 ), 
        .B0(n2659), .B1(\addr_calc/fft_read_calc/count[22] ), .Y(n1012) );
  XNOR2X4TS U2590 ( .A(\DP_OP_159_297_3515/n913 ), .B(n1678), .Y(n1702) );
  AO22X4TS U2591 ( .A0(n1759), .A1(\addr_calc/fir_write_calc/counter/N61 ), 
        .B0(n1266), .B1(\addr_calc/fir_write_calc/count[18] ), .Y(n1112) );
  BUFX4TS U2592 ( .A(n2654), .Y(n2649) );
  XNOR2X4TS U2593 ( .A(\DP_OP_159_297_3515/n948 ), .B(
        \DP_OP_159_297_3515/n862 ), .Y(n1703) );
  AND2X8TS U2594 ( .A(\DP_OP_158_296_6262/n62 ), .B(\DP_OP_158_296_6262/n3 ), 
        .Y(n1715) );
  BUFX6TS U2595 ( .A(n2794), .Y(n2661) );
  XNOR2X4TS U2596 ( .A(n1731), .B(n2558), .Y(\DP_OP_158_296_6262/n133 ) );
  OR4X6TS U2597 ( .A(n783), .B(n2793), .C(\data_cntl/N63 ), .D(n2588), .Y(
        n1704) );
  NOR2X2TS U2598 ( .A(\DP_OP_159_297_3515/n714 ), .B(\DP_OP_159_297_3515/n723 ), .Y(\DP_OP_159_297_3515/n712 ) );
  CLKINVX3TS U2599 ( .A(n2787), .Y(n1705) );
  CLKINVX3TS U2600 ( .A(n2787), .Y(n1706) );
  INVX2TS U2601 ( .A(n1458), .Y(n1707) );
  INVX2TS U2602 ( .A(n1705), .Y(n1708) );
  INVX2TS U2603 ( .A(n1458), .Y(n1709) );
  INVX2TS U2604 ( .A(n1706), .Y(n1710) );
  INVX2TS U2605 ( .A(n1705), .Y(n1711) );
  INVX2TS U2606 ( .A(n1706), .Y(n1712) );
  INVX2TS U2607 ( .A(n1458), .Y(n1713) );
  INVX2TS U2608 ( .A(n1705), .Y(n1714) );
  NAND2X8TS U2609 ( .A(n1715), .B(n1716), .Y(
        \addr_calc/fir_read_calc/counter/N38 ) );
  AND2X8TS U2610 ( .A(\DP_OP_158_296_6262/n179 ), .B(\DP_OP_158_296_6262/n280 ), .Y(n1716) );
  NAND2X2TS U2611 ( .A(\DP_OP_159_297_3515/n907 ), .B(n1791), .Y(
        \DP_OP_159_297_3515/n906 ) );
  XOR2X4TS U2612 ( .A(\DP_OP_159_297_3515/n1010 ), .B(n1682), .Y(n2618) );
  NOR2X2TS U2613 ( .A(n1717), .B(\DP_OP_158_296_6262/n1834 ), .Y(
        \DP_OP_158_296_6262/n1833 ) );
  NAND2X2TS U2614 ( .A(n1788), .B(\DP_OP_159_297_3515/n997 ), .Y(
        \DP_OP_159_297_3515/n996 ) );
  OR2X8TS U2615 ( .A(\DP_OP_158_296_6262/n2011 ), .B(
        \DP_OP_158_296_6262/n1987 ), .Y(n1728) );
  AO22X4TS U2616 ( .A0(n1762), .A1(\addr_calc/fir_write_calc/counter/N62 ), 
        .B0(n1267), .B1(n1670), .Y(n1111) );
  AO22X4TS U2617 ( .A0(n1723), .A1(\addr_calc/fft_write_calc/counter/N53 ), 
        .B0(n2666), .B1(n1932), .Y(n1056) );
  AO22X4TS U2618 ( .A0(n1722), .A1(\addr_calc/fft_write_calc/counter/N52 ), 
        .B0(n2664), .B1(n1934), .Y(n1057) );
  AO22X4TS U2619 ( .A0(n1725), .A1(\addr_calc/fft_write_calc/counter/N50 ), 
        .B0(n2667), .B1(n1936), .Y(n1059) );
  AO22X4TS U2620 ( .A0(n1725), .A1(\addr_calc/fft_write_calc/counter/N58 ), 
        .B0(n2667), .B1(n1976), .Y(n1051) );
  XNOR2X4TS U2621 ( .A(\DP_OP_158_296_6262/n1881 ), .B(n2344), .Y(n1731) );
  INVX3TS U2622 ( .A(n1820), .Y(n1826) );
  AO22X4TS U2623 ( .A0(n1723), .A1(\addr_calc/fft_write_calc/counter/N64 ), 
        .B0(n2668), .B1(\addr_calc/fft_write_calc/count[21] ), .Y(n1045) );
  AO22X4TS U2624 ( .A0(n1727), .A1(\addr_calc/fft_write_calc/counter/N62 ), 
        .B0(n2664), .B1(\addr_calc/fft_write_calc/count[19] ), .Y(n1047) );
  XNOR2X4TS U2625 ( .A(\DP_OP_159_297_3515/n996 ), .B(
        \DP_OP_159_297_3515/n869 ), .Y(n2616) );
  NAND2X2TS U2626 ( .A(n1787), .B(\DP_OP_159_297_3515/n1004 ), .Y(
        \DP_OP_159_297_3515/n1003 ) );
  INVX2TS U2627 ( .A(n1819), .Y(n1822) );
  INVX2TS U2628 ( .A(n1819), .Y(n1823) );
  INVX2TS U2629 ( .A(n1819), .Y(n1821) );
  AO22X4TS U2630 ( .A0(n1145), .A1(\addr_calc/fft_write_calc/counter/N56 ), 
        .B0(n2665), .B1(n1927), .Y(n1053) );
  AO22X4TS U2631 ( .A0(n1725), .A1(\addr_calc/fft_write_calc/counter/N55 ), 
        .B0(n2665), .B1(n2023), .Y(n1054) );
  INVX2TS U2632 ( .A(n1765), .Y(n1770) );
  BUFX6TS U2633 ( .A(n2812), .Y(n2680) );
  AO22X4TS U2634 ( .A0(n1151), .A1(\addr_calc/fir_read_calc/counter/N65 ), 
        .B0(n1744), .B1(\addr_calc/fir_read_calc/count[22] ), .Y(n1076) );
  XOR2X4TS U2635 ( .A(\DP_OP_158_296_6262/n1847 ), .B(n2330), .Y(n1775) );
  MXI2X2TS U2636 ( .A(n2806), .B(\addr_calc/fir_write_calc/counter/N43 ), .S0(
        n1265), .Y(n1130) );
  NOR2X2TS U2637 ( .A(n1781), .B(n1737), .Y(n2787) );
  XNOR2X4TS U2638 ( .A(n1697), .B(n2048), .Y(\DP_OP_159_297_3515/n593 ) );
  NAND2X2TS U2639 ( .A(n1787), .B(\DP_OP_159_297_3515/n1018 ), .Y(
        \DP_OP_159_297_3515/n1017 ) );
  NOR2X4TS U2640 ( .A(\DP_OP_159_297_3515/n610 ), .B(\DP_OP_159_297_3515/n593 ), .Y(\DP_OP_159_297_3515/n591 ) );
  NOR2X4TS U2641 ( .A(\DP_OP_158_296_6262/n104 ), .B(\DP_OP_158_296_6262/n119 ), .Y(\DP_OP_158_296_6262/n102 ) );
  INVX2TS U2642 ( .A(n1757), .Y(n1759) );
  NAND2X2TS U2643 ( .A(n1788), .B(\DP_OP_159_297_3515/n990 ), .Y(
        \DP_OP_159_297_3515/n989 ) );
  NOR2X2TS U2644 ( .A(\DP_OP_158_296_6262/n255 ), .B(\DP_OP_158_296_6262/n242 ), .Y(\DP_OP_158_296_6262/n240 ) );
  BUFX6TS U2645 ( .A(n2654), .Y(n2652) );
  AO22X4TS U2646 ( .A0(n1708), .A1(\addr_calc/iir_read_calc/counter/N62 ), 
        .B0(n2651), .B1(n2556), .Y(n952) );
  NOR2X2TS U2647 ( .A(\addr_calc/iir_read_calc/count[12] ), .B(n2410), .Y(
        \add_x_19_4/n131 ) );
  INVX2TS U2648 ( .A(n1766), .Y(n1771) );
  INVX4TS U2649 ( .A(n2813), .Y(n1766) );
  BUFX4TS U2650 ( .A(n2794), .Y(n2660) );
  AO22X4TS U2651 ( .A0(n1767), .A1(\addr_calc/iir_write_calc/counter/N51 ), 
        .B0(n2680), .B1(n2041), .Y(n994) );
  AO22X4TS U2652 ( .A0(n1711), .A1(\addr_calc/iir_read_calc/counter/N54 ), 
        .B0(n2649), .B1(\addr_calc/iir_read_calc/count[11] ), .Y(n960) );
  AO22X4TS U2653 ( .A0(n1774), .A1(\addr_calc/iir_write_calc/counter/N52 ), 
        .B0(n2673), .B1(n2562), .Y(n993) );
  BUFX6TS U2654 ( .A(n2679), .Y(n2675) );
  CLKINVX6TS U2655 ( .A(n2807), .Y(n1819) );
  AO22X4TS U2656 ( .A0(n1710), .A1(\addr_calc/iir_read_calc/counter/N63 ), 
        .B0(n2651), .B1(\addr_calc/iir_read_calc/count[20] ), .Y(n951) );
  AO22X4TS U2657 ( .A0(n1825), .A1(\addr_calc/fir_read_calc/counter/N66 ), 
        .B0(n1744), .B1(n2558), .Y(n1075) );
  XNOR2X4TS U2658 ( .A(\DP_OP_158_296_6262/n1826 ), .B(n2325), .Y(n1778) );
  NOR2X2TS U2659 ( .A(n1796), .B(\DP_OP_158_296_6262/n1827 ), .Y(
        \DP_OP_158_296_6262/n1826 ) );
  XNOR2X4TS U2660 ( .A(\DP_OP_158_296_6262/n1957 ), .B(n2368), .Y(n1756) );
  NOR2X2TS U2661 ( .A(n1693), .B(n1455), .Y(\DP_OP_158_296_6262/n1957 ) );
  INVX2TS U2662 ( .A(\add_x_22_4/n74 ), .Y(n1785) );
  NAND2X2TS U2663 ( .A(\addr_calc/iir_read_calc/count[12] ), .B(n2410), .Y(
        \add_x_19_4/n132 ) );
  XNOR2X4TS U2664 ( .A(\DP_OP_158_296_6262/n833 ), .B(n2582), .Y(
        \DP_OP_158_296_6262/n87 ) );
  NOR2X4TS U2665 ( .A(\DP_OP_158_296_6262/n181 ), .B(\DP_OP_158_296_6262/n238 ), .Y(\DP_OP_158_296_6262/n179 ) );
  NAND2X2TS U2666 ( .A(\DP_OP_158_296_6262/n264 ), .B(
        \DP_OP_158_296_6262/n240 ), .Y(\DP_OP_158_296_6262/n238 ) );
  NAND2X4TS U2667 ( .A(\DP_OP_158_296_6262/n183 ), .B(
        \DP_OP_158_296_6262/n215 ), .Y(\DP_OP_158_296_6262/n181 ) );
  NOR2X4TS U2668 ( .A(\DP_OP_158_296_6262/n202 ), .B(\DP_OP_158_296_6262/n185 ), .Y(\DP_OP_158_296_6262/n183 ) );
  BUFX8TS U2669 ( .A(n2812), .Y(n2679) );
  INVX6TS U2670 ( .A(\DP_OP_158_296_6262/n2051 ), .Y(\DP_OP_158_296_6262/n838 ) );
  XNOR2X2TS U2671 ( .A(n1729), .B(n1884), .Y(\DP_OP_158_296_6262/n217 ) );
  AO22X4TS U2672 ( .A0(n1694), .A1(\addr_calc/fft_write_calc/counter/N51 ), 
        .B0(n2664), .B1(n2026), .Y(n1058) );
  AO22X4TS U2673 ( .A0(n1721), .A1(\addr_calc/fft_write_calc/counter/N66 ), 
        .B0(n2666), .B1(n2555), .Y(n1043) );
  AO22X4TS U2674 ( .A0(n1725), .A1(\addr_calc/fft_write_calc/counter/N71 ), 
        .B0(n2669), .B1(n2557), .Y(n1038) );
  BUFX6TS U2675 ( .A(n2671), .Y(n2669) );
  AO22X4TS U2676 ( .A0(n1694), .A1(\addr_calc/fft_write_calc/counter/N46 ), 
        .B0(n2663), .B1(n2568), .Y(n1063) );
  BUFX6TS U2677 ( .A(n2671), .Y(n2663) );
  BUFX4TS U2678 ( .A(n2671), .Y(n2665) );
  XNOR2X4TS U2679 ( .A(n2619), .B(n2044), .Y(\DP_OP_159_297_3515/n694 ) );
  XNOR2X4TS U2680 ( .A(\DP_OP_159_297_3515/n1017 ), .B(
        \DP_OP_158_296_6262/n1952 ), .Y(n2619) );
  NAND2X2TS U2681 ( .A(\DP_OP_158_296_6262/n37 ), .B(n1653), .Y(
        \DP_OP_158_296_6262/n18 ) );
  XNOR2X2TS U2682 ( .A(n1655), .B(\addr_calc/fir_read_calc/count[25] ), .Y(
        \DP_OP_158_296_6262/n104 ) );
  XNOR2X4TS U2683 ( .A(n1718), .B(n1983), .Y(\DP_OP_158_296_6262/n119 ) );
  AND4X1TS U2684 ( .A(\add_x_22_4/n57 ), .B(\add_x_22_4/n64 ), .C(
        \add_x_22_4/n67 ), .D(\add_x_22_4/n71 ), .Y(n817) );
  INVX2TS U2685 ( .A(\addr_calc/iir_read_calc/count[15] ), .Y(\add_x_22_4/n64 ) );
  NAND2X2TS U2686 ( .A(\DP_OP_159_297_3515/n921 ), .B(n1791), .Y(
        \DP_OP_159_297_3515/n920 ) );
  XNOR2X2TS U2687 ( .A(n1654), .B(n1881), .Y(\DP_OP_158_296_6262/n185 ) );
  XOR2X4TS U2688 ( .A(\DP_OP_158_296_6262/n2004 ), .B(n1493), .Y(n2595) );
  XNOR2X4TS U2689 ( .A(\add_x_19_4/n57 ), .B(\add_x_19_4/n5 ), .Y(
        \addr_calc/iir_read_addr[27] ) );
  XOR2X4TS U2690 ( .A(\DP_OP_158_296_6262/n1833 ), .B(n2341), .Y(
        \DP_OP_158_296_6262/n2060 ) );
  NOR2X2TS U2691 ( .A(\DP_OP_158_296_6262/n217 ), .B(\DP_OP_158_296_6262/n230 ), .Y(\DP_OP_158_296_6262/n215 ) );
  AO22X4TS U2692 ( .A0(n1708), .A1(\addr_calc/iir_read_calc/counter/N55 ), 
        .B0(n2648), .B1(n1785), .Y(n959) );
  AO22X4TS U2693 ( .A0(n1712), .A1(\addr_calc/iir_read_calc/counter/N57 ), 
        .B0(n2648), .B1(n1784), .Y(n957) );
  NOR2X2TS U2694 ( .A(\DP_OP_158_296_6262/n1998 ), .B(n2366), .Y(
        \DP_OP_158_296_6262/n1991 ) );
  NAND2X2TS U2695 ( .A(\DP_OP_159_297_3515/n956 ), .B(
        \DP_OP_159_297_3515/n930 ), .Y(\DP_OP_159_297_3515/n852 ) );
  NOR2X4TS U2696 ( .A(n1794), .B(\DP_OP_158_296_6262/n1917 ), .Y(
        \DP_OP_158_296_6262/n1916 ) );
  NAND2X2TS U2697 ( .A(\DP_OP_158_296_6262/n66 ), .B(\DP_OP_158_296_6262/n102 ), .Y(\DP_OP_158_296_6262/n64 ) );
  NAND2X2TS U2698 ( .A(\DP_OP_158_296_6262/n159 ), .B(
        \DP_OP_158_296_6262/n131 ), .Y(\DP_OP_158_296_6262/n129 ) );
  BUFX6TS U2699 ( .A(n2654), .Y(n2647) );
  NOR2X4TS U2700 ( .A(n1794), .B(\DP_OP_158_296_6262/n1910 ), .Y(
        \DP_OP_158_296_6262/n1909 ) );
  NOR2X2TS U2701 ( .A(n1728), .B(\DP_OP_158_296_6262/n1944 ), .Y(
        \DP_OP_158_296_6262/n1943 ) );
  XOR2X4TS U2702 ( .A(\DP_OP_158_296_6262/n1895 ), .B(n1679), .Y(
        \DP_OP_158_296_6262/n2051 ) );
  AOI21X4TS U2703 ( .A0(\addr_calc/fir_read_calc/counter/N38 ), .A1(
        data_to_fir), .B0(n2060), .Y(n2809) );
  XOR2X4TS U2704 ( .A(\DP_OP_158_296_6262/n1916 ), .B(n1523), .Y(
        \DP_OP_158_296_6262/n2048 ) );
  INVX2TS U2705 ( .A(n1812), .Y(n1813) );
  INVX2TS U2706 ( .A(n1806), .Y(n1807) );
  NAND2X2TS U2707 ( .A(\DP_OP_159_297_3515/n692 ), .B(
        \DP_OP_159_297_3515/n712 ), .Y(\DP_OP_159_297_3515/n690 ) );
  NOR2X2TS U2708 ( .A(\DP_OP_159_297_3515/n705 ), .B(\DP_OP_159_297_3515/n694 ), .Y(\DP_OP_159_297_3515/n692 ) );
  XNOR2X4TS U2709 ( .A(\DP_OP_159_297_3515/n1031 ), .B(
        \DP_OP_158_296_6262/n1966 ), .Y(n2621) );
  AO22X4TS U2710 ( .A0(n1773), .A1(\addr_calc/iir_write_calc/counter/N65 ), 
        .B0(n2674), .B1(n2579), .Y(n980) );
  AO22X4TS U2711 ( .A0(n1824), .A1(\addr_calc/fir_read_calc/counter/N71 ), 
        .B0(n1460), .B1(\addr_calc/fir_read_calc/count[28] ), .Y(n1070) );
  MXI2X2TS U2712 ( .A(n2792), .B(n2791), .S0(n2672), .Y(n1002) );
  XOR2X4TS U2713 ( .A(\DP_OP_159_297_3515/n976 ), .B(
        \DP_OP_158_296_6262/n1911 ), .Y(\DP_OP_159_297_3515/n1128 ) );
  BUFX4TS U2714 ( .A(\DP_OP_159_297_3515/n1039 ), .Y(n1786) );
  MXI2X2TS U2715 ( .A(n2811), .B(n2810), .S0(n1674), .Y(n1098) );
  AO22X4TS U2716 ( .A0(n1753), .A1(\addr_calc/fft_read_calc/counter/N73 ), 
        .B0(n1476), .B1(\addr_calc/fft_read_calc/count[30] ), .Y(n1004) );
  CLKINVX3TS U2717 ( .A(n1782), .Y(n1790) );
  INVX2TS U2718 ( .A(n2419), .Y(n2420) );
  INVXLTS U2719 ( .A(instruction[26]), .Y(n1798) );
  INVXLTS U2720 ( .A(instruction[27]), .Y(n1800) );
  INVXLTS U2721 ( .A(instruction[15]), .Y(n1802) );
  INVXLTS U2722 ( .A(instruction[28]), .Y(n1804) );
  INVXLTS U2723 ( .A(filesize[28]), .Y(n1806) );
  INVXLTS U2724 ( .A(filesize[29]), .Y(n1808) );
  INVXLTS U2725 ( .A(offset[9]), .Y(n1810) );
  INVXLTS U2726 ( .A(n1810), .Y(n1811) );
  INVXLTS U2727 ( .A(offset[8]), .Y(n2471) );
  INVXLTS U2728 ( .A(filesize[17]), .Y(n1812) );
  INVXLTS U2729 ( .A(filesize[24]), .Y(n1814) );
  INVXLTS U2730 ( .A(filesize[27]), .Y(n1816) );
  NAND2X1TS U2731 ( .A(n1813), .B(n1523), .Y(\DP_OP_159_297_3515/n971 ) );
  INVXLTS U2732 ( .A(n1531), .Y(\DP_OP_159_297_3515/n964 ) );
  AO21X1TS U2733 ( .A0(\add_x_19_5/n179 ), .A1(\add_x_19_5/n187 ), .B0(
        \add_x_19_5/n180 ), .Y(n1818) );
  AO22X4TS U2734 ( .A0(n1727), .A1(\addr_calc/fft_write_calc/counter/N73 ), 
        .B0(n2669), .B1(\addr_calc/fft_write_calc/count[30] ), .Y(n1036) );
  AO22X4TS U2735 ( .A0(n1823), .A1(\addr_calc/fir_read_calc/counter/N72 ), 
        .B0(n1747), .B1(\addr_calc/fir_read_calc/count[29] ), .Y(n1069) );
  INVX2TS U2736 ( .A(\DP_OP_159_297_3515/n956 ), .Y(\DP_OP_159_297_3515/n957 )
         );
  AO22X4TS U2737 ( .A0(n1824), .A1(\addr_calc/fir_read_calc/counter/N57 ), 
        .B0(n1744), .B1(\addr_calc/fir_read_calc/count[14] ), .Y(n1084) );
  NAND2X2TS U2738 ( .A(\DP_OP_159_297_3515/n956 ), .B(
        \DP_OP_159_297_3515/n930 ), .Y(n2551) );
  NOR2X2TS U2739 ( .A(\DP_OP_159_297_3515/n943 ), .B(\DP_OP_159_297_3515/n931 ), .Y(\DP_OP_159_297_3515/n930 ) );
  AO22X4TS U2740 ( .A0(n1707), .A1(\addr_calc/iir_read_calc/counter/N61 ), 
        .B0(n2651), .B1(\addr_calc/iir_read_calc/count[18] ), .Y(n953) );
  NOR2X1TS U2741 ( .A(\addr_calc/fft_read_calc/count[6] ), .B(n2428), .Y(
        \add_x_19_0/n165 ) );
  NOR2X1TS U2742 ( .A(\addr_calc/iir_read_calc/count[23] ), .B(n2468), .Y(
        \add_x_19_4/n78 ) );
  CLKBUFX2TS U2743 ( .A(\addr_calc/fir_write_calc/count[30] ), .Y(n1836) );
  INVX2TS U2744 ( .A(\addr_calc/iir_read_calc/count[30] ), .Y(n1843) );
  INVX2TS U2745 ( .A(\addr_calc/iir_read_calc/count[31] ), .Y(n1846) );
  INVX2TS U2746 ( .A(n1846), .Y(n1847) );
  INVX2TS U2747 ( .A(n1848), .Y(n1849) );
  CLKBUFX2TS U2748 ( .A(\addr_calc/iir_write_calc/count[30] ), .Y(n1854) );
  CLKBUFX2TS U2749 ( .A(\addr_calc/iir_write_calc/count[31] ), .Y(n1857) );
  INVX2TS U2750 ( .A(n1858), .Y(n1859) );
  INVX2TS U2751 ( .A(n2815), .Y(n1860) );
  INVX2TS U2752 ( .A(\addr_calc/fir_write_calc/count[3] ), .Y(
        \add_x_22_3/n114 ) );
  CLKBUFX2TS U2753 ( .A(\addr_calc/fir_write_calc/count[1] ), .Y(n1868) );
  NOR2X1TS U2754 ( .A(\addr_calc/fir_read_calc/count[27] ), .B(n2499), .Y(
        \add_x_19_2/n55 ) );
  INVX2TS U2755 ( .A(\addr_calc/fir_write_calc/count[10] ), .Y(
        \add_x_22_3/n84 ) );
  INVX2TS U2756 ( .A(\addr_calc/fir_read_calc/count[25] ), .Y(n1875) );
  INVX2TS U2757 ( .A(n1875), .Y(n1876) );
  INVX2TS U2758 ( .A(\addr_calc/fir_write_calc/count[15] ), .Y(n1882) );
  INVX2TS U2759 ( .A(\addr_calc/fir_write_calc/count[17] ), .Y(n1885) );
  INVX2TS U2760 ( .A(n1885), .Y(n1886) );
  INVX2TS U2761 ( .A(\addr_calc/fir_read_calc/count[16] ), .Y(n1887) );
  NOR4XLTS U2762 ( .A(\addr_calc/fir_write_calc/count[30] ), .B(
        \addr_calc/fir_write_calc/count[2] ), .C(n1833), .D(
        \addr_calc/fir_write_calc/count[28] ), .Y(n864) );
  INVX2TS U2763 ( .A(\add_x_22_4/n121 ), .Y(n1898) );
  INVX2TS U2764 ( .A(\addr_calc/iir_read_calc/count[1] ), .Y(\add_x_22_4/n121 ) );
  CLKBUFX2TS U2765 ( .A(\addr_calc/iir_read_calc/count[4] ), .Y(n1903) );
  INVX2TS U2766 ( .A(\addr_calc/fft_write_calc/count[27] ), .Y(n1912) );
  INVX2TS U2767 ( .A(n1912), .Y(n1913) );
  INVX2TS U2768 ( .A(\addr_calc/fft_write_calc/count[25] ), .Y(n1914) );
  INVX2TS U2769 ( .A(n1914), .Y(n1915) );
  INVX2TS U2770 ( .A(\addr_calc/fft_write_calc/count[21] ), .Y(n1917) );
  INVX2TS U2771 ( .A(n1921), .Y(n1922) );
  INVX2TS U2772 ( .A(n1925), .Y(n1926) );
  INVX2TS U2773 ( .A(n1928), .Y(n1929) );
  INVX2TS U2774 ( .A(\add_x_22_5/n121 ), .Y(n1931) );
  INVX2TS U2775 ( .A(\addr_calc/iir_write_calc/count[4] ), .Y(
        \add_x_22_5/n109 ) );
  INVX2TS U2776 ( .A(\add_x_22_1/n109 ), .Y(n1939) );
  AO22X4TS U2777 ( .A0(n1722), .A1(\addr_calc/fft_write_calc/counter/N47 ), 
        .B0(n2663), .B1(n1939), .Y(n1062) );
  INVX2TS U2778 ( .A(\addr_calc/fft_write_calc/count[4] ), .Y(
        \add_x_22_1/n109 ) );
  INVX2TS U2779 ( .A(\add_x_22_1/n121 ), .Y(n1941) );
  INVX2TS U2780 ( .A(\addr_calc/fft_write_calc/count[1] ), .Y(
        \add_x_22_1/n121 ) );
  INVX2TS U2781 ( .A(\addr_calc/fft_read_calc/count[25] ), .Y(n1946) );
  INVX2TS U2782 ( .A(\addr_calc/fft_read_calc/count[23] ), .Y(n1949) );
  INVX2TS U2783 ( .A(n1949), .Y(n1950) );
  INVX2TS U2784 ( .A(\addr_calc/fft_read_calc/count[19] ), .Y(n1955) );
  INVX2TS U2785 ( .A(n1957), .Y(n1958) );
  INVX2TS U2786 ( .A(\addr_calc/fft_read_calc/count[17] ), .Y(n1959) );
  INVX2TS U2787 ( .A(\addr_calc/iir_write_calc/count[21] ), .Y(n1961) );
  INVX2TS U2788 ( .A(n1961), .Y(n1962) );
  INVX2TS U2789 ( .A(\addr_calc/fft_read_calc/count[15] ), .Y(n1963) );
  INVX2TS U2790 ( .A(n1964), .Y(n1965) );
  INVX2TS U2791 ( .A(\addr_calc/fft_read_calc/count[13] ), .Y(n1966) );
  INVX2TS U2792 ( .A(n1966), .Y(n1967) );
  INVX2TS U2793 ( .A(\addr_calc/iir_write_calc/count[25] ), .Y(n1968) );
  INVX2TS U2794 ( .A(\addr_calc/fft_read_calc/count[7] ), .Y(n1975) );
  CLKBUFX2TS U2795 ( .A(\addr_calc/fft_read_calc/count[5] ), .Y(n1977) );
  INVX2TS U2796 ( .A(\add_x_22_0/n114 ), .Y(n1978) );
  INVX2TS U2797 ( .A(\add_x_22_0/n121 ), .Y(n1979) );
  INVX2TS U2798 ( .A(\addr_calc/fft_read_calc/count[1] ), .Y(\add_x_22_0/n121 ) );
  INVX2TS U2799 ( .A(n2494), .Y(n1980) );
  NOR2X1TS U2800 ( .A(\addr_calc/fft_write_calc/count[9] ), .B(n2495), .Y(
        \add_x_19_1/n151 ) );
  INVX2TS U2801 ( .A(n1811), .Y(n2494) );
  CLKBUFX2TS U2802 ( .A(\addr_calc/fir_write_calc/count[0] ), .Y(n1986) );
  INVX2TS U2803 ( .A(\addr_calc/fir_read_calc/count[18] ), .Y(n1987) );
  INVX2TS U2804 ( .A(n1987), .Y(n1988) );
  INVX2TS U2805 ( .A(\addr_calc/fir_read_calc/count[14] ), .Y(n1991) );
  CLKBUFX2TS U2806 ( .A(\addr_calc/fir_write_calc/count[6] ), .Y(n1993) );
  CLKBUFX2TS U2807 ( .A(\addr_calc/fir_write_calc/count[8] ), .Y(n1996) );
  INVX2TS U2808 ( .A(\addr_calc/fir_write_calc/count[12] ), .Y(n1998) );
  INVX2TS U2809 ( .A(\addr_calc/fir_read_calc/count[6] ), .Y(\add_x_22_2/n101 ) );
  INVX2TS U2810 ( .A(n2002), .Y(n2003) );
  INVX2TS U2811 ( .A(\add_x_22_2/n117 ), .Y(n2004) );
  INVX2TS U2812 ( .A(\addr_calc/fir_read_calc/count[2] ), .Y(\add_x_22_2/n117 ) );
  INVX2TS U2813 ( .A(\addr_calc/fir_read_calc/count[0] ), .Y(n2810) );
  INVX2TS U2814 ( .A(\addr_calc/fir_write_calc/count[20] ), .Y(n2008) );
  INVX2TS U2815 ( .A(\addr_calc/fft_write_calc/count[24] ), .Y(n2010) );
  INVX2TS U2816 ( .A(n2010), .Y(n2011) );
  INVX2TS U2817 ( .A(\addr_calc/fir_write_calc/count[22] ), .Y(n2012) );
  INVX2TS U2818 ( .A(\addr_calc/fft_write_calc/count[22] ), .Y(n2013) );
  INVX2TS U2819 ( .A(\add_x_22_4/n117 ), .Y(n2015) );
  INVX2TS U2820 ( .A(\addr_calc/iir_read_calc/count[2] ), .Y(\add_x_22_4/n117 ) );
  INVX2TS U2821 ( .A(\addr_calc/fft_write_calc/count[20] ), .Y(n2016) );
  INVX2TS U2822 ( .A(\addr_calc/iir_read_calc/count[6] ), .Y(\add_x_22_4/n101 ) );
  INVX2TS U2823 ( .A(\addr_calc/fft_write_calc/count[18] ), .Y(n2019) );
  CLKBUFX2TS U2824 ( .A(\addr_calc/fft_write_calc/count[14] ), .Y(n2022) );
  AO22X4TS U2825 ( .A0(n1723), .A1(\addr_calc/fft_write_calc/counter/N57 ), 
        .B0(n2665), .B1(n2022), .Y(n1052) );
  NAND2X1TS U2826 ( .A(\addr_calc/fft_write_calc/count[8] ), .B(n2472), .Y(
        \add_x_19_1/n155 ) );
  INVX2TS U2827 ( .A(\addr_calc/iir_read_calc/count[20] ), .Y(n2027) );
  INVX2TS U2828 ( .A(n2029), .Y(n2030) );
  NOR2X1TS U2829 ( .A(\addr_calc/iir_read_calc/count[22] ), .B(n2464), .Y(
        \add_x_19_4/n81 ) );
  INVX2TS U2830 ( .A(\add_x_22_1/n117 ), .Y(n2032) );
  INVX2TS U2831 ( .A(\addr_calc/fft_write_calc/count[2] ), .Y(
        \add_x_22_1/n117 ) );
  INVX2TS U2832 ( .A(\addr_calc/iir_read_calc/count[24] ), .Y(n2033) );
  INVX2TS U2833 ( .A(n2033), .Y(n2034) );
  INVX2TS U2834 ( .A(\add_x_22_5/n117 ), .Y(n2036) );
  INVX2TS U2835 ( .A(\addr_calc/iir_write_calc/count[2] ), .Y(
        \add_x_22_5/n117 ) );
  INVX2TS U2836 ( .A(\addr_calc/fft_read_calc/count[24] ), .Y(n2037) );
  INVX2TS U2837 ( .A(n2037), .Y(n2038) );
  INVX2TS U2838 ( .A(\addr_calc/iir_write_calc/count[6] ), .Y(
        \add_x_22_5/n101 ) );
  INVX2TS U2839 ( .A(\addr_calc/fft_read_calc/count[14] ), .Y(n2042) );
  INVX2TS U2840 ( .A(\addr_calc/iir_write_calc/count[12] ), .Y(
        \add_x_22_5/n74 ) );
  INVX2TS U2841 ( .A(\addr_calc/fft_read_calc/count[12] ), .Y(n2045) );
  INVX2TS U2842 ( .A(n2050), .Y(n2051) );
  INVX2TS U2843 ( .A(\addr_calc/fft_read_calc/count[6] ), .Y(\add_x_22_0/n101 ) );
  INVX2TS U2844 ( .A(\add_x_22_0/n117 ), .Y(n2056) );
  INVX2TS U2845 ( .A(\addr_calc/fft_read_calc/count[2] ), .Y(\add_x_22_0/n117 ) );
  INVX2TS U2846 ( .A(n1783), .Y(\DP_OP_158_296_6262/n1875 ) );
  INVXLTS U2847 ( .A(n2066), .Y(n2059) );
  INVXLTS U2848 ( .A(n2062), .Y(iir_enable) );
  INVXLTS U2849 ( .A(n2065), .Y(n2067) );
  INVXLTS U2850 ( .A(n2070), .Y(n2071) );
  INVXLTS U2851 ( .A(n2070), .Y(n2073) );
  INVXLTS U2852 ( .A(instruction[12]), .Y(n2075) );
  INVXLTS U2853 ( .A(instruction[17]), .Y(n2077) );
  INVXLTS U2854 ( .A(instruction[13]), .Y(n2079) );
  INVXLTS U2855 ( .A(instruction[22]), .Y(n2081) );
  INVXLTS U2856 ( .A(instruction[6]), .Y(n2083) );
  INVXLTS U2857 ( .A(instruction[23]), .Y(n2085) );
  INVXLTS U2858 ( .A(instruction[10]), .Y(n2087) );
  INVXLTS U2859 ( .A(instruction[11]), .Y(n2089) );
  INVXLTS U2860 ( .A(instruction[7]), .Y(n2091) );
  INVXLTS U2861 ( .A(instruction[18]), .Y(n2093) );
  INVXLTS U2862 ( .A(instruction[4]), .Y(n2094) );
  INVXLTS U2863 ( .A(instruction[20]), .Y(n2096) );
  INVXLTS U2864 ( .A(instruction[16]), .Y(n2098) );
  INVXLTS U2865 ( .A(instruction[21]), .Y(n2100) );
  INVXLTS U2866 ( .A(instruction[3]), .Y(n2102) );
  INVXLTS U2867 ( .A(instruction[25]), .Y(n2104) );
  INVXLTS U2868 ( .A(instruction[14]), .Y(n2106) );
  INVXLTS U2869 ( .A(instruction[19]), .Y(n2108) );
  INVXLTS U2870 ( .A(instruction[8]), .Y(n2109) );
  INVXLTS U2871 ( .A(instruction[24]), .Y(n2111) );
  INVXLTS U2872 ( .A(instruction[5]), .Y(n2113) );
  INVXLTS U2873 ( .A(reset), .Y(n2115) );
  INVXLTS U2874 ( .A(fir_data_in[15]), .Y(n2117) );
  INVXLTS U2875 ( .A(fir_data_in[16]), .Y(n2119) );
  INVXLTS U2876 ( .A(fir_data_in[14]), .Y(n2121) );
  INVXLTS U2877 ( .A(fir_data_in[17]), .Y(n2123) );
  INVXLTS U2878 ( .A(fir_data_in[13]), .Y(n2125) );
  INVXLTS U2879 ( .A(fir_data_in[18]), .Y(n2127) );
  INVXLTS U2880 ( .A(fir_data_in[12]), .Y(n2129) );
  INVXLTS U2881 ( .A(fir_data_in[19]), .Y(n2131) );
  INVXLTS U2882 ( .A(fir_data_in[11]), .Y(n2133) );
  INVXLTS U2883 ( .A(fir_data_in[20]), .Y(n2135) );
  INVXLTS U2884 ( .A(fir_data_in[10]), .Y(n2137) );
  INVXLTS U2885 ( .A(fir_data_in[21]), .Y(n2139) );
  INVXLTS U2886 ( .A(fir_data_in[9]), .Y(n2141) );
  INVXLTS U2887 ( .A(fir_data_in[22]), .Y(n2143) );
  INVXLTS U2888 ( .A(fir_data_in[8]), .Y(n2145) );
  INVXLTS U2889 ( .A(fir_data_in[23]), .Y(n2147) );
  INVXLTS U2890 ( .A(fir_data_in[7]), .Y(n2149) );
  INVXLTS U2891 ( .A(fir_data_in[24]), .Y(n2151) );
  INVXLTS U2892 ( .A(fir_data_in[6]), .Y(n2153) );
  INVXLTS U2893 ( .A(fir_data_in[25]), .Y(n2155) );
  INVXLTS U2894 ( .A(fir_data_in[5]), .Y(n2157) );
  INVXLTS U2895 ( .A(fir_data_in[26]), .Y(n2159) );
  INVXLTS U2896 ( .A(fir_data_in[4]), .Y(n2161) );
  INVXLTS U2897 ( .A(fir_data_in[27]), .Y(n2163) );
  INVXLTS U2898 ( .A(fir_data_in[3]), .Y(n2165) );
  INVXLTS U2899 ( .A(fir_data_in[28]), .Y(n2167) );
  INVXLTS U2900 ( .A(fir_data_in[2]), .Y(n2169) );
  INVXLTS U2901 ( .A(fir_data_in[29]), .Y(n2171) );
  INVXLTS U2902 ( .A(fir_data_in[1]), .Y(n2173) );
  INVXLTS U2903 ( .A(fir_data_in[30]), .Y(n2175) );
  INVXLTS U2904 ( .A(fir_data_in[0]), .Y(n2177) );
  INVXLTS U2905 ( .A(fir_data_in[31]), .Y(n2179) );
  INVXLTS U2906 ( .A(iir_data_in[31]), .Y(n2181) );
  INVXLTS U2907 ( .A(fft_data_in[0]), .Y(n2183) );
  INVXLTS U2908 ( .A(iir_data_in[30]), .Y(n2185) );
  INVXLTS U2909 ( .A(fft_data_in[1]), .Y(n2187) );
  INVXLTS U2910 ( .A(iir_data_in[29]), .Y(n2189) );
  INVXLTS U2911 ( .A(fft_data_in[2]), .Y(n2191) );
  INVXLTS U2912 ( .A(iir_data_in[28]), .Y(n2193) );
  INVXLTS U2913 ( .A(fft_data_in[3]), .Y(n2195) );
  INVXLTS U2914 ( .A(iir_data_in[27]), .Y(n2197) );
  INVXLTS U2915 ( .A(fft_data_in[4]), .Y(n2199) );
  INVXLTS U2916 ( .A(iir_data_in[26]), .Y(n2201) );
  INVXLTS U2917 ( .A(fft_data_in[5]), .Y(n2203) );
  INVXLTS U2918 ( .A(iir_data_in[25]), .Y(n2205) );
  INVXLTS U2919 ( .A(fft_data_in[6]), .Y(n2207) );
  INVXLTS U2920 ( .A(iir_data_in[24]), .Y(n2209) );
  INVXLTS U2921 ( .A(fft_data_in[7]), .Y(n2211) );
  INVXLTS U2922 ( .A(iir_data_in[23]), .Y(n2213) );
  INVXLTS U2923 ( .A(fft_data_in[8]), .Y(n2215) );
  INVXLTS U2924 ( .A(iir_data_in[22]), .Y(n2217) );
  INVXLTS U2925 ( .A(fft_data_in[9]), .Y(n2219) );
  INVXLTS U2926 ( .A(iir_data_in[21]), .Y(n2221) );
  INVXLTS U2927 ( .A(fft_data_in[10]), .Y(n2223) );
  INVXLTS U2928 ( .A(iir_data_in[20]), .Y(n2225) );
  INVXLTS U2929 ( .A(fft_data_in[11]), .Y(n2227) );
  INVXLTS U2930 ( .A(iir_data_in[19]), .Y(n2229) );
  INVXLTS U2931 ( .A(fft_data_in[12]), .Y(n2231) );
  INVXLTS U2932 ( .A(iir_data_in[18]), .Y(n2233) );
  INVXLTS U2933 ( .A(fft_data_in[13]), .Y(n2235) );
  INVXLTS U2934 ( .A(iir_data_in[17]), .Y(n2237) );
  INVXLTS U2935 ( .A(fft_data_in[14]), .Y(n2239) );
  INVXLTS U2936 ( .A(iir_data_in[16]), .Y(n2241) );
  INVXLTS U2937 ( .A(fft_data_in[15]), .Y(n2243) );
  INVXLTS U2938 ( .A(iir_data_in[15]), .Y(n2245) );
  INVXLTS U2939 ( .A(fft_data_in[16]), .Y(n2247) );
  INVXLTS U2940 ( .A(iir_data_in[14]), .Y(n2249) );
  INVXLTS U2941 ( .A(fft_data_in[17]), .Y(n2251) );
  INVXLTS U2942 ( .A(iir_data_in[13]), .Y(n2253) );
  INVXLTS U2943 ( .A(fft_data_in[18]), .Y(n2255) );
  INVXLTS U2944 ( .A(iir_data_in[12]), .Y(n2257) );
  INVXLTS U2945 ( .A(fft_data_in[19]), .Y(n2259) );
  INVXLTS U2946 ( .A(iir_data_in[11]), .Y(n2261) );
  INVXLTS U2947 ( .A(fft_data_in[20]), .Y(n2263) );
  INVXLTS U2948 ( .A(iir_data_in[10]), .Y(n2265) );
  INVXLTS U2949 ( .A(fft_data_in[21]), .Y(n2267) );
  INVXLTS U2950 ( .A(iir_data_in[9]), .Y(n2269) );
  INVXLTS U2951 ( .A(fft_data_in[22]), .Y(n2271) );
  INVXLTS U2952 ( .A(iir_data_in[8]), .Y(n2273) );
  INVXLTS U2953 ( .A(fft_data_in[23]), .Y(n2275) );
  INVXLTS U2954 ( .A(iir_data_in[7]), .Y(n2277) );
  INVXLTS U2955 ( .A(fft_data_in[24]), .Y(n2279) );
  INVXLTS U2956 ( .A(iir_data_in[6]), .Y(n2281) );
  INVXLTS U2957 ( .A(fft_data_in[25]), .Y(n2283) );
  INVXLTS U2958 ( .A(iir_data_in[5]), .Y(n2285) );
  INVXLTS U2959 ( .A(fft_data_in[26]), .Y(n2287) );
  INVXLTS U2960 ( .A(iir_data_in[4]), .Y(n2289) );
  INVXLTS U2961 ( .A(fft_data_in[27]), .Y(n2291) );
  INVXLTS U2962 ( .A(iir_data_in[3]), .Y(n2293) );
  INVXLTS U2963 ( .A(fft_data_in[28]), .Y(n2295) );
  INVXLTS U2964 ( .A(iir_data_in[2]), .Y(n2297) );
  INVXLTS U2965 ( .A(fft_data_in[29]), .Y(n2299) );
  INVXLTS U2966 ( .A(iir_data_in[1]), .Y(n2301) );
  INVXLTS U2967 ( .A(fft_data_in[30]), .Y(n2303) );
  INVXLTS U2968 ( .A(iir_data_in[0]), .Y(n2305) );
  INVXLTS U2969 ( .A(fft_data_in[31]), .Y(n2307) );
  INVX2TS U2970 ( .A(\DP_OP_158_296_6262/n1830 ), .Y(n2341) );
  INVXLTS U2971 ( .A(instruction[0]), .Y(n2309) );
  INVXLTS U2972 ( .A(instruction[1]), .Y(n2311) );
  INVXLTS U2973 ( .A(to_fir_full), .Y(n2312) );
  INVXLTS U2974 ( .A(from_fir_full), .Y(n2314) );
  INVXLTS U2975 ( .A(from_fft_empty), .Y(n2316) );
  INVXLTS U2976 ( .A(to_fft_full), .Y(n2318) );
  INVXLTS U2977 ( .A(to_fft_empty), .Y(n2320) );
  INVXLTS U2978 ( .A(to_iir_full), .Y(n2322) );
  INVXLTS U2979 ( .A(filesize[31]), .Y(n2324) );
  INVXLTS U2980 ( .A(from_iir_full), .Y(n2326) );
  INVXLTS U2981 ( .A(from_fir_empty), .Y(n2328) );
  INVXLTS U2982 ( .A(to_fir_empty), .Y(n2331) );
  INVXLTS U2983 ( .A(from_fft_full), .Y(n2333) );
  INVXLTS U2984 ( .A(instruction[2]), .Y(n2335) );
  INVXLTS U2985 ( .A(from_iir_empty), .Y(n2337) );
  INVXLTS U2986 ( .A(to_iir_empty), .Y(n2339) );
  INVXLTS U2987 ( .A(filesize[30]), .Y(\DP_OP_158_296_6262/n1830 ) );
  INVX2TS U2988 ( .A(n1808), .Y(n2342) );
  INVXLTS U2989 ( .A(data_bus[15]), .Y(n2345) );
  INVXLTS U2990 ( .A(data_bus[19]), .Y(n2347) );
  INVXLTS U2991 ( .A(data_bus[11]), .Y(n2349) );
  INVXLTS U2992 ( .A(data_bus[23]), .Y(n2351) );
  INVXLTS U2993 ( .A(data_bus[7]), .Y(n2353) );
  INVXLTS U2994 ( .A(data_bus[27]), .Y(n2355) );
  INVXLTS U2995 ( .A(data_bus[3]), .Y(n2357) );
  INVXLTS U2996 ( .A(data_bus[31]), .Y(n2359) );
  INVXLTS U2997 ( .A(n1487), .Y(\DP_OP_159_297_3515/n873 ) );
  INVXLTS U2998 ( .A(n1493), .Y(\DP_OP_159_297_3515/n879 ) );
  INVXLTS U2999 ( .A(n1529), .Y(\DP_OP_159_297_3515/n868 ) );
  INVXLTS U3000 ( .A(n1489), .Y(\DP_OP_159_297_3515/n877 ) );
  NOR2XLTS U3001 ( .A(\DP_OP_159_297_3515/n1074 ), .B(n2363), .Y(
        \DP_OP_159_297_3515/n1069 ) );
  INVXLTS U3002 ( .A(n1813), .Y(\DP_OP_159_297_3515/n867 ) );
  INVXLTS U3003 ( .A(n1525), .Y(\DP_OP_159_297_3515/n815 ) );
  INVXLTS U3004 ( .A(filesize[1]), .Y(n2373) );
  INVX2TS U3005 ( .A(n2373), .Y(n2374) );
  INVXLTS U3006 ( .A(offset[26]), .Y(n2375) );
  INVXLTS U3007 ( .A(offset[31]), .Y(n2379) );
  INVXLTS U3008 ( .A(offset[28]), .Y(n2383) );
  INVXLTS U3009 ( .A(offset[29]), .Y(n2387) );
  INVXLTS U3010 ( .A(offset[0]), .Y(n2391) );
  INVXLTS U3011 ( .A(offset[4]), .Y(n2395) );
  INVXLTS U3012 ( .A(offset[16]), .Y(n2399) );
  INVXLTS U3013 ( .A(offset[11]), .Y(n2403) );
  INVXLTS U3014 ( .A(offset[12]), .Y(n2407) );
  INVXLTS U3015 ( .A(offset[10]), .Y(n2411) );
  INVXLTS U3016 ( .A(offset[13]), .Y(n2415) );
  INVXLTS U3017 ( .A(offset[7]), .Y(n2419) );
  INVXLTS U3018 ( .A(offset[14]), .Y(n2423) );
  INVXLTS U3019 ( .A(offset[6]), .Y(n2427) );
  INVXLTS U3020 ( .A(offset[18]), .Y(n2431) );
  INVXLTS U3021 ( .A(offset[3]), .Y(n2435) );
  INVXLTS U3022 ( .A(offset[20]), .Y(n2439) );
  INVXLTS U3023 ( .A(offset[2]), .Y(n2443) );
  INVXLTS U3024 ( .A(offset[21]), .Y(n2447) );
  INVXLTS U3025 ( .A(offset[1]), .Y(n2451) );
  INVXLTS U3026 ( .A(n2451), .Y(n2452) );
  INVXLTS U3027 ( .A(offset[30]), .Y(n2455) );
  INVXLTS U3028 ( .A(offset[24]), .Y(n2459) );
  INVXLTS U3029 ( .A(offset[22]), .Y(n2463) );
  INVXLTS U3030 ( .A(offset[23]), .Y(n2467) );
  INVXLTS U3031 ( .A(offset[15]), .Y(n2474) );
  INVXLTS U3032 ( .A(offset[17]), .Y(n2478) );
  INVXLTS U3033 ( .A(offset[5]), .Y(n2482) );
  INVXLTS U3034 ( .A(offset[19]), .Y(n2486) );
  INVXLTS U3035 ( .A(offset[25]), .Y(n2490) );
  INVX2TS U3036 ( .A(n2494), .Y(n2495) );
  INVX2TS U3037 ( .A(n2494), .Y(n2496) );
  INVXLTS U3038 ( .A(offset[27]), .Y(n2497) );
  INVXLTS U3039 ( .A(data_bus[30]), .Y(n2501) );
  INVXLTS U3040 ( .A(data_bus[26]), .Y(n2503) );
  INVXLTS U3041 ( .A(data_bus[22]), .Y(n2505) );
  INVXLTS U3042 ( .A(data_bus[18]), .Y(n2507) );
  INVXLTS U3043 ( .A(data_bus[14]), .Y(n2509) );
  INVXLTS U3044 ( .A(data_bus[10]), .Y(n2511) );
  INVXLTS U3045 ( .A(data_bus[6]), .Y(n2513) );
  INVXLTS U3046 ( .A(data_bus[2]), .Y(n2515) );
  INVXLTS U3047 ( .A(data_bus[29]), .Y(n2517) );
  INVXLTS U3048 ( .A(data_bus[25]), .Y(n2519) );
  INVXLTS U3049 ( .A(data_bus[21]), .Y(n2521) );
  INVXLTS U3050 ( .A(data_bus[17]), .Y(n2523) );
  INVXLTS U3051 ( .A(data_bus[13]), .Y(n2525) );
  INVXLTS U3052 ( .A(data_bus[9]), .Y(n2527) );
  INVXLTS U3053 ( .A(data_bus[5]), .Y(n2529) );
  INVXLTS U3054 ( .A(data_bus[1]), .Y(n2531) );
  INVXLTS U3055 ( .A(data_bus[28]), .Y(n2533) );
  INVXLTS U3056 ( .A(data_bus[24]), .Y(n2535) );
  INVXLTS U3057 ( .A(data_bus[20]), .Y(n2537) );
  INVXLTS U3058 ( .A(data_bus[16]), .Y(n2539) );
  INVXLTS U3059 ( .A(data_bus[12]), .Y(n2541) );
  INVXLTS U3060 ( .A(data_bus[8]), .Y(n2543) );
  INVXLTS U3061 ( .A(data_bus[4]), .Y(n2545) );
  INVXLTS U3062 ( .A(data_bus[0]), .Y(n2547) );
  CLKBUFX2TS U3063 ( .A(\addr_calc/fir_read_calc/count[31] ), .Y(n2549) );
  CLKBUFX2TS U3064 ( .A(\addr_calc/fir_write_calc/count[31] ), .Y(n2550) );
  NOR2XLTS U3065 ( .A(\addr_calc/fft_read_calc/count[4] ), .B(n2396), .Y(
        \add_x_19_0/n175 ) );
  INVX2TS U3066 ( .A(\add_x_22_0/n57 ), .Y(n2554) );
  NOR2XLTS U3067 ( .A(\addr_calc/fft_read_calc/count[16] ), .B(n2402), .Y(
        \add_x_19_0/n110 ) );
  INVX2TS U3068 ( .A(\add_x_22_1/n30 ), .Y(n2555) );
  INVX2TS U3069 ( .A(\add_x_22_4/n46 ), .Y(n2556) );
  INVX2TS U3070 ( .A(\add_x_22_1/n7 ), .Y(n2557) );
  INVX2TS U3071 ( .A(\add_x_22_2/n30 ), .Y(n2558) );
  NOR2X1TS U3072 ( .A(\addr_calc/fir_read_calc/count[23] ), .B(n2468), .Y(
        \add_x_19_2/n78 ) );
  INVX2TS U3073 ( .A(\add_x_22_0/n7 ), .Y(n2559) );
  INVX2TS U3074 ( .A(\add_x_22_0/n89 ), .Y(n2560) );
  INVX2TS U3075 ( .A(\add_x_22_4/n7 ), .Y(n2561) );
  INVX2TS U3076 ( .A(\add_x_22_5/n89 ), .Y(n2562) );
  INVX2TS U3077 ( .A(\add_x_22_3/n30 ), .Y(n2563) );
  INVX2TS U3078 ( .A(\add_x_22_3/n57 ), .Y(n2564) );
  NAND2X1TS U3079 ( .A(\addr_calc/fir_write_calc/count[16] ), .B(n2402), .Y(
        \add_x_19_3/n111 ) );
  INVX2TS U3080 ( .A(\add_x_22_4/n30 ), .Y(n2565) );
  INVX2TS U3081 ( .A(\add_x_22_1/n57 ), .Y(n2567) );
  NAND2X1TS U3082 ( .A(\addr_calc/fft_write_calc/count[16] ), .B(n2402), .Y(
        \add_x_19_1/n111 ) );
  INVX2TS U3083 ( .A(\add_x_22_1/n114 ), .Y(n2568) );
  INVX2TS U3084 ( .A(\add_x_22_5/n67 ), .Y(n2570) );
  INVX2TS U3085 ( .A(\add_x_22_5/n49 ), .Y(n2571) );
  INVX2TS U3086 ( .A(\add_x_22_0/n40 ), .Y(n2572) );
  INVX2TS U3087 ( .A(\add_x_22_5/n15 ), .Y(n2573) );
  INVX2TS U3088 ( .A(\add_x_22_1/n15 ), .Y(n2574) );
  INVX2TS U3089 ( .A(\add_x_22_0/n15 ), .Y(n2575) );
  INVX2TS U3090 ( .A(\add_x_22_4/n15 ), .Y(n2576) );
  INVX2TS U3091 ( .A(\add_x_22_3/n22 ), .Y(n2577) );
  INVX2TS U3092 ( .A(n2791), .Y(n2578) );
  XNOR2X1TS U3093 ( .A(\addr_calc/iir_write_calc/count[0] ), .B(
        \DP_OP_159_297_3515/n815 ), .Y(\DP_OP_159_297_3515/n778 ) );
  INVX2TS U3094 ( .A(\add_x_22_5/n33 ), .Y(n2579) );
  INVX2TS U3095 ( .A(n2786), .Y(n2580) );
  INVX2TS U3096 ( .A(\add_x_22_3/n15 ), .Y(n2581) );
  NOR4XLTS U3097 ( .A(\addr_calc/fir_write_calc/count[25] ), .B(
        \addr_calc/fir_write_calc/count[26] ), .C(n1835), .D(
        \addr_calc/fir_write_calc/count[24] ), .Y(n863) );
  INVX2TS U3098 ( .A(\add_x_22_2/n15 ), .Y(n2582) );
  NOR2X1TS U3099 ( .A(\addr_calc/fir_read_calc/count[26] ), .B(n2376), .Y(
        \add_x_19_2/n58 ) );
  INVX2TS U3100 ( .A(\add_x_22_4/n92 ), .Y(n2583) );
  INVX2TS U3101 ( .A(n2584), .Y(n2587) );
  INVX2TS U3102 ( .A(n2584), .Y(n2586) );
  AOI211XLTS U3103 ( .A0(n2321), .A1(n938), .B0(n2317), .C0(n2587), .Y(
        \data_cntl/N252 ) );
  INVX2TS U3104 ( .A(\addr_calc/fft_read_calc/count[16] ), .Y(\add_x_22_0/n57 ) );
  INVX2TS U3105 ( .A(\add_x_22_0/n24 ), .Y(\add_x_22_0/n23 ) );
  XNOR2X1TS U3106 ( .A(\add_x_22_2/n121 ), .B(n2007), .Y(
        \addr_calc/fir_read_calc/counter/N44 ) );
  INVX2TS U3107 ( .A(\addr_calc/fir_read_calc/count[27] ), .Y(\add_x_22_2/n12 ) );
  INVX2TS U3108 ( .A(\addr_calc/fir_read_calc/count[23] ), .Y(\add_x_22_2/n30 ) );
  INVX2TS U3109 ( .A(\addr_calc/fir_read_calc/count[26] ), .Y(\add_x_22_2/n15 ) );
  INVX2TS U3110 ( .A(\addr_calc/fir_write_calc/count[16] ), .Y(
        \add_x_22_3/n57 ) );
  INVX2TS U3111 ( .A(\addr_calc/fir_write_calc/count[24] ), .Y(
        \add_x_22_3/n22 ) );
  INVX2TS U3112 ( .A(\addr_calc/iir_write_calc/count[17] ), .Y(
        \add_x_22_5/n53 ) );
  INVX2TS U3113 ( .A(\addr_calc/iir_write_calc/count[22] ), .Y(
        \add_x_22_5/n33 ) );
  INVX2TS U3114 ( .A(\addr_calc/fft_write_calc/count[16] ), .Y(
        \add_x_22_1/n57 ) );
  INVX2TS U3115 ( .A(\addr_calc/iir_read_calc/count[22] ), .Y(\add_x_22_4/n33 ) );
  INVX2TS U3116 ( .A(\addr_calc/iir_read_calc/count[16] ), .Y(\add_x_22_4/n57 ) );
  INVXLTS U3117 ( .A(\addr_calc/iir_read_calc/count[5] ), .Y(\add_x_22_4/n105 ) );
  XNOR2X1TS U3118 ( .A(n2372), .B(\addr_calc/fir_read_calc/count[0] ), .Y(
        \DP_OP_158_296_6262/n375 ) );
  XOR2X1TS U3119 ( .A(n2596), .B(n2004), .Y(n2590) );
  XOR2X1TS U3120 ( .A(n2593), .B(\addr_calc/fir_read_calc/count[6] ), .Y(n2591) );
  XOR2X1TS U3121 ( .A(n2599), .B(n1908), .Y(n2592) );
  XOR2X1TS U3122 ( .A(\DP_OP_158_296_6262/n855 ), .B(
        \addr_calc/fir_read_calc/count[4] ), .Y(n2600) );
  XOR2X1TS U3123 ( .A(n2595), .B(n1904), .Y(n2601) );
  INVXLTS U3124 ( .A(n1138), .Y(\DP_OP_158_296_6262/n1972 ) );
  XOR2X1TS U3125 ( .A(n2374), .B(n1648), .Y(n2597) );
  INVX2TS U3126 ( .A(\DP_OP_158_296_6262/n2011 ), .Y(
        \DP_OP_158_296_6262/n2010 ) );
  INVX2TS U3127 ( .A(\DP_OP_158_296_6262/n2034 ), .Y(\DP_OP_158_296_6262/n855 ) );
  INVXLTS U3128 ( .A(\DP_OP_158_296_6262/n1862 ), .Y(
        \DP_OP_158_296_6262/n1863 ) );
  INVXLTS U3129 ( .A(\DP_OP_158_296_6262/n1918 ), .Y(
        \DP_OP_158_296_6262/n1917 ) );
  INVX2TS U3130 ( .A(n1797), .Y(\DP_OP_158_296_6262/n2020 ) );
  INVX2TS U3131 ( .A(\DP_OP_158_296_6262/n1903 ), .Y(
        \DP_OP_158_296_6262/n1904 ) );
  INVX2TS U3132 ( .A(\DP_OP_158_296_6262/n1792 ), .Y(
        \DP_OP_158_296_6262/n1849 ) );
  XOR2X4TS U3133 ( .A(\DP_OP_158_296_6262/n1874 ), .B(n1815), .Y(
        \DP_OP_158_296_6262/n2054 ) );
  NOR2X2TS U3134 ( .A(\DP_OP_158_296_6262/n68 ), .B(\DP_OP_158_296_6262/n87 ), 
        .Y(\DP_OP_158_296_6262/n66 ) );
  NOR2X2TS U3135 ( .A(\DP_OP_158_296_6262/n18 ), .B(\DP_OP_158_296_6262/n5 ), 
        .Y(\DP_OP_158_296_6262/n3 ) );
  NOR2X2TS U3136 ( .A(\DP_OP_158_296_6262/n54 ), .B(\DP_OP_158_296_6262/n39 ), 
        .Y(\DP_OP_158_296_6262/n37 ) );
  NOR2X2TS U3137 ( .A(\DP_OP_158_296_6262/n174 ), .B(\DP_OP_158_296_6262/n161 ), .Y(\DP_OP_158_296_6262/n159 ) );
  NAND2X1TS U3138 ( .A(\DP_OP_159_297_3515/n893 ), .B(n1789), .Y(
        \DP_OP_159_297_3515/n892 ) );
  XOR2X1TS U3139 ( .A(n2612), .B(\addr_calc/iir_write_calc/count[2] ), .Y(
        n2604) );
  XOR2X1TS U3140 ( .A(n2610), .B(n2039), .Y(n2605) );
  XOR2X1TS U3141 ( .A(n2624), .B(n1935), .Y(n2606) );
  XOR2X1TS U3142 ( .A(\DP_OP_159_297_3515/n1051 ), .B(
        \DP_OP_159_297_3515/n877 ), .Y(n2609) );
  XOR2X1TS U3143 ( .A(\DP_OP_159_297_3515/n1074 ), .B(n2363), .Y(n2611) );
  XOR2X1TS U3144 ( .A(n1680), .B(n2374), .Y(n2612) );
  XNOR2X1TS U3145 ( .A(\DP_OP_159_297_3515/n1063 ), .B(
        \DP_OP_159_297_3515/n879 ), .Y(n2623) );
  XNOR2X1TS U3146 ( .A(\DP_OP_159_297_3515/n1069 ), .B(
        \DP_OP_159_297_3515/n880 ), .Y(n2624) );
  XOR2X1TS U3147 ( .A(n2623), .B(n1686), .Y(n2626) );
  INVX2TS U3148 ( .A(\DP_OP_159_297_3515/n1011 ), .Y(
        \DP_OP_159_297_3515/n1012 ) );
  INVX2TS U3149 ( .A(\DP_OP_159_297_3515/n1064 ), .Y(
        \DP_OP_159_297_3515/n1063 ) );
  INVXLTS U3150 ( .A(n1650), .Y(\DP_OP_159_297_3515/n1074 ) );
  INVXLTS U3151 ( .A(\DP_OP_159_297_3515/n915 ), .Y(\DP_OP_159_297_3515/n916 )
         );
  INVXLTS U3152 ( .A(\DP_OP_159_297_3515/n998 ), .Y(\DP_OP_159_297_3515/n999 )
         );
  XOR2X4TS U3153 ( .A(\DP_OP_159_297_3515/n906 ), .B(n2330), .Y(
        \DP_OP_159_297_3515/n1138 ) );
  NOR2X2TS U3154 ( .A(\DP_OP_159_297_3515/n742 ), .B(\DP_OP_159_297_3515/n758 ), .Y(\DP_OP_159_297_3515/n740 ) );
  NAND2X2TS U3155 ( .A(\DP_OP_159_297_3515/n728 ), .B(
        \DP_OP_159_297_3515/n740 ), .Y(\DP_OP_159_297_3515/n726 ) );
  XNOR2X4TS U3156 ( .A(n1662), .B(\addr_calc/iir_write_calc/count[19] ), .Y(
        \DP_OP_159_297_3515/n610 ) );
  OR2X2TS U3157 ( .A(\addr_calc/fft_read_calc/count[29] ), .B(n2389), .Y(n2628) );
  OR2X2TS U3158 ( .A(n1856), .B(n2382), .Y(n2627) );
  INVX2TS U3159 ( .A(\add_x_19_0/n69 ), .Y(\add_x_19_0/n68 ) );
  XNOR2X4TS U3160 ( .A(\add_x_19_0/n35 ), .B(\add_x_19_0/n1 ), .Y(
        \addr_calc/fft_read_addr[31] ) );
  OAI21X2TS U3161 ( .A0(\add_x_19_0/n38 ), .A1(\add_x_19_0/n36 ), .B0(
        \add_x_19_0/n37 ), .Y(\add_x_19_0/n35 ) );
  NAND2X2TS U3162 ( .A(n2058), .B(n2394), .Y(\add_x_19_0/n191 ) );
  INVX2TS U3163 ( .A(\add_x_19_5/n157 ), .Y(\add_x_19_5/n156 ) );
  OR2X2TS U3164 ( .A(n1851), .B(n2389), .Y(n2629) );
  INVX2TS U3165 ( .A(\add_x_19_5/n113 ), .Y(\add_x_19_5/n112 ) );
  INVX2TS U3166 ( .A(\add_x_19_5/n92 ), .Y(\add_x_19_5/n91 ) );
  INVX2TS U3167 ( .A(\add_x_19_5/n69 ), .Y(\add_x_19_5/n68 ) );
  OAI21X1TS U3168 ( .A0(\add_x_19_5/n105 ), .A1(\add_x_19_5/n111 ), .B0(
        \add_x_19_5/n106 ), .Y(\add_x_19_5/n104 ) );
  OAI21X2TS U3169 ( .A0(\add_x_19_5/n113 ), .A1(\add_x_19_5/n70 ), .B0(
        \add_x_19_5/n71 ), .Y(\add_x_19_5/n69 ) );
  INVX2TS U3170 ( .A(\add_x_19_3/n157 ), .Y(\add_x_19_3/n156 ) );
  OR2X2TS U3171 ( .A(n1833), .B(n2390), .Y(n2631) );
  OAI21X2TS U3172 ( .A0(\add_x_19_3/n38 ), .A1(\add_x_19_3/n36 ), .B0(
        \add_x_19_3/n37 ), .Y(\add_x_19_3/n35 ) );
  AOI21X1TS U3173 ( .A0(\add_x_19_3/n69 ), .A1(\add_x_19_3/n61 ), .B0(
        \add_x_19_3/n62 ), .Y(\add_x_19_3/n60 ) );
  INVXLTS U3174 ( .A(\add_x_19_1/n139 ), .Y(\add_x_19_1/n212 ) );
  OR2X2TS U3175 ( .A(\addr_calc/fft_write_calc/count[29] ), .B(n2388), .Y(
        n2632) );
  OR2X2TS U3176 ( .A(n1842), .B(n2390), .Y(n2633) );
  INVX2TS U3177 ( .A(\add_x_19_2/n69 ), .Y(\add_x_19_2/n68 ) );
  INVX2TS U3178 ( .A(\add_x_19_4/n157 ), .Y(\add_x_19_4/n156 ) );
  OR2X2TS U3179 ( .A(\addr_calc/iir_read_calc/count[29] ), .B(n2389), .Y(n2634) );
  INVX2TS U3180 ( .A(\add_x_19_4/n134 ), .Y(\add_x_19_4/n133 ) );
  INVXLTS U3181 ( .A(\add_x_19_4/n178 ), .Y(\add_x_19_4/n177 ) );
  AO22X4TS U3182 ( .A0(n1710), .A1(\addr_calc/iir_read_calc/counter/N74 ), 
        .B0(n2652), .B1(\addr_calc/iir_read_calc/count[31] ), .Y(n972) );
  AO22X4TS U3183 ( .A0(n1774), .A1(\addr_calc/iir_write_calc/counter/N57 ), 
        .B0(n2675), .B1(n2570), .Y(n988) );
  AO22X4TS U3184 ( .A0(n1714), .A1(\addr_calc/iir_read_calc/counter/N73 ), 
        .B0(n2650), .B1(n1684), .Y(n941) );
  AO22X4TS U3185 ( .A0(n1767), .A1(\addr_calc/iir_write_calc/counter/N50 ), 
        .B0(n2674), .B1(n1683), .Y(n995) );
  AO22X4TS U3186 ( .A0(n1768), .A1(\addr_calc/iir_write_calc/counter/N55 ), 
        .B0(n2674), .B1(n2044), .Y(n990) );
  AO22X4TS U3187 ( .A0(n1770), .A1(\addr_calc/iir_write_calc/counter/N53 ), 
        .B0(n2673), .B1(n1940), .Y(n992) );
  AO22X4TS U3188 ( .A0(n1771), .A1(\addr_calc/iir_write_calc/counter/N72 ), 
        .B0(n2676), .B1(n1851), .Y(n973) );
  AO22X4TS U3189 ( .A0(n1711), .A1(\addr_calc/iir_read_calc/counter/N53 ), 
        .B0(n2648), .B1(n1909), .Y(n961) );
  AO22X4TS U3190 ( .A0(n1709), .A1(\addr_calc/iir_read_calc/counter/N51 ), 
        .B0(n2649), .B1(n2583), .Y(n963) );
  AO22X4TS U3191 ( .A0(n1711), .A1(\addr_calc/iir_read_calc/counter/N52 ), 
        .B0(n2649), .B1(n1685), .Y(n962) );
  CLKINVX6TS U3192 ( .A(n1649), .Y(n787) );
  CLKINVX6TS U3193 ( .A(\addr_calc/fir_write_calc/counter/N38 ), .Y(n785) );
  AO22X4TS U3194 ( .A0(n1713), .A1(\addr_calc/iir_read_calc/counter/N58 ), 
        .B0(n2650), .B1(n2566), .Y(n956) );
  NOR4XLTS U3195 ( .A(\addr_calc/fir_read_calc/count[27] ), .B(
        \addr_calc/fir_read_calc/count[26] ), .C(n1876), .D(n1983), .Y(n878)
         );
  NOR4XLTS U3196 ( .A(\addr_calc/fir_read_calc/count[5] ), .B(n1906), .C(n1908), .D(\addr_calc/fir_read_calc/count[31] ), .Y(n876) );
  NOR4XLTS U3197 ( .A(n1867), .B(\addr_calc/fir_write_calc/count[4] ), .C(
        n1866), .D(\addr_calc/fir_write_calc/count[31] ), .Y(n861) );
  NOR4XLTS U3198 ( .A(n1859), .B(n2056), .C(n1863), .D(
        \addr_calc/fft_read_calc/count[28] ), .Y(n831) );
  NOR4XLTS U3199 ( .A(\addr_calc/fft_read_calc/count[27] ), .B(
        \addr_calc/fft_read_calc/count[26] ), .C(
        \addr_calc/fft_read_calc/count[25] ), .D(n2038), .Y(n830) );
  NOR4XLTS U3200 ( .A(n1977), .B(n2552), .C(n1978), .D(n1856), .Y(n828) );
  NOR4XLTS U3201 ( .A(n1849), .B(n2032), .C(n1853), .D(
        \addr_calc/fft_write_calc/count[28] ), .Y(n845) );
  NOR4XLTS U3202 ( .A(\addr_calc/fft_write_calc/count[27] ), .B(
        \addr_calc/fft_write_calc/count[26] ), .C(
        \addr_calc/fft_write_calc/count[25] ), .D(
        \addr_calc/fft_write_calc/count[24] ), .Y(n844) );
  NOR4XLTS U3203 ( .A(n1479), .B(n1939), .C(n2568), .D(n1845), .Y(n842) );
  NOR4XLTS U3204 ( .A(\addr_calc/iir_write_calc/count[27] ), .B(
        \addr_calc/iir_write_calc/count[26] ), .C(
        \addr_calc/iir_write_calc/count[25] ), .D(
        \addr_calc/iir_write_calc/count[24] ), .Y(n917) );
  BUFX3TS U3205 ( .A(n2654), .Y(n2653) );
  NOR4XLTS U3206 ( .A(\addr_calc/iir_read_calc/count[30] ), .B(n2015), .C(
        n1840), .D(\addr_calc/iir_read_calc/count[28] ), .Y(n813) );
  NOR4XLTS U3207 ( .A(\addr_calc/iir_read_calc/count[27] ), .B(
        \addr_calc/iir_read_calc/count[26] ), .C(
        \addr_calc/iir_read_calc/count[25] ), .D(n2034), .Y(n812) );
  BUFX3TS U3208 ( .A(n2670), .Y(n2667) );
  NOR4XLTS U3209 ( .A(n2553), .B(n1903), .C(\addr_calc/iir_read_calc/count[3] ), .D(n1847), .Y(n810) );
  NOR4XLTS U3210 ( .A(\addr_calc/iir_write_calc/count[5] ), .B(n1935), .C(
        \addr_calc/iir_write_calc/count[3] ), .D(
        \addr_calc/iir_write_calc/count[31] ), .Y(n915) );
  NOR2X1TS U3211 ( .A(n2800), .B(n2799), .Y(n2808) );
  NOR2X1TS U3212 ( .A(n2802), .B(n2801), .Y(n2804) );
  NOR2X1TS U3213 ( .A(n2784), .B(n2783), .Y(n2785) );
  BUFX3TS U3214 ( .A(n2661), .Y(n2657) );
  BUFX3TS U3215 ( .A(n2670), .Y(n2664) );
  BUFX3TS U3216 ( .A(n2670), .Y(n2666) );
  AO22X2TS U3217 ( .A0(n1151), .A1(\addr_calc/fir_read_calc/counter/N62 ), 
        .B0(n1671), .B1(n1881), .Y(n1079) );
  AO22X2TS U3218 ( .A0(n1762), .A1(\addr_calc/fir_write_calc/counter/N72 ), 
        .B0(n1260), .B1(\addr_calc/fir_write_calc/count[29] ), .Y(n1101) );
  AO22X2TS U3219 ( .A0(n1755), .A1(\addr_calc/fft_read_calc/counter/N58 ), 
        .B0(n2658), .B1(n1689), .Y(n1019) );
  AO22X2TS U3220 ( .A0(n1755), .A1(\addr_calc/fft_read_calc/counter/N72 ), 
        .B0(n2658), .B1(n1863), .Y(n1005) );
  AO22X2TS U3221 ( .A0(n1726), .A1(\addr_calc/fft_write_calc/counter/N72 ), 
        .B0(n2669), .B1(n1853), .Y(n1037) );
  CLKBUFX2TS U3222 ( .A(n2725), .Y(n2719) );
  CLKBUFX2TS U3223 ( .A(n2725), .Y(n2720) );
  CLKBUFX2TS U3224 ( .A(n2725), .Y(n2724) );
  CLKBUFX2TS U3225 ( .A(n451), .Y(n2725) );
  INVXLTS U3226 ( .A(\data_cntl/N159 ), .Y(n451) );
  CLKBUFX2TS U3227 ( .A(n323), .Y(n2739) );
  CLKBUFX2TS U3228 ( .A(n323), .Y(n2741) );
  CLKBUFX2TS U3229 ( .A(n259), .Y(n2747) );
  CLKBUFX2TS U3230 ( .A(n259), .Y(n2749) );
  CLKBUFX2TS U3231 ( .A(n195), .Y(n2755) );
  CLKBUFX2TS U3232 ( .A(n195), .Y(n2757) );
  CLKBUFX2TS U3233 ( .A(n131), .Y(n2762) );
  CLKBUFX2TS U3234 ( .A(n131), .Y(n2763) );
  CLKBUFX2TS U3235 ( .A(n2698), .Y(n2692) );
  CLKBUFX2TS U3236 ( .A(n2698), .Y(n2693) );
  CLKBUFX2TS U3237 ( .A(n2698), .Y(n2696) );
  CLKBUFX2TS U3238 ( .A(n2698), .Y(n2697) );
  CLKBUFX2TS U3239 ( .A(n643), .Y(n2698) );
  INVXLTS U3240 ( .A(\data_cntl/N63 ), .Y(n643) );
  CLKBUFX2TS U3241 ( .A(n2716), .Y(n2710) );
  CLKBUFX2TS U3242 ( .A(n2716), .Y(n2711) );
  CLKBUFX2TS U3243 ( .A(n2716), .Y(n2714) );
  CLKBUFX2TS U3244 ( .A(n2716), .Y(n2715) );
  CLKBUFX2TS U3245 ( .A(n515), .Y(n2716) );
  INVXLTS U3246 ( .A(\data_cntl/N99 ), .Y(n515) );
  CLKBUFX2TS U3247 ( .A(n2734), .Y(n2728) );
  CLKBUFX2TS U3248 ( .A(n2734), .Y(n2729) );
  CLKBUFX2TS U3249 ( .A(n2734), .Y(n2732) );
  CLKBUFX2TS U3250 ( .A(n2734), .Y(n2733) );
  CLKBUFX2TS U3251 ( .A(n387), .Y(n2734) );
  INVXLTS U3252 ( .A(\data_cntl/N191 ), .Y(n387) );
  CLKBUFX2TS U3253 ( .A(n2689), .Y(n2683) );
  CLKBUFX2TS U3254 ( .A(n2689), .Y(n2684) );
  CLKBUFX2TS U3255 ( .A(n2689), .Y(n2688) );
  CLKBUFX2TS U3256 ( .A(n707), .Y(n2689) );
  INVXLTS U3257 ( .A(\data_cntl/N9 ), .Y(n707) );
  CLKBUFX2TS U3258 ( .A(n2707), .Y(n2701) );
  CLKBUFX2TS U3259 ( .A(n2707), .Y(n2702) );
  CLKBUFX2TS U3260 ( .A(n2707), .Y(n2706) );
  CLKBUFX2TS U3261 ( .A(n579), .Y(n2707) );
  INVXLTS U3262 ( .A(\data_cntl/N95 ), .Y(n579) );
  CLKBUFX2TS U3263 ( .A(n195), .Y(n2753) );
  CLKBUFX2TS U3264 ( .A(n131), .Y(n2765) );
  CLKBUFX2TS U3265 ( .A(n131), .Y(n2761) );
  INVXLTS U3266 ( .A(\addr_calc/N99 ), .Y(n131) );
  CLKBUFX2TS U3267 ( .A(n67), .Y(n2770) );
  CLKBUFX2TS U3268 ( .A(n323), .Y(n2738) );
  CLKBUFX2TS U3269 ( .A(n259), .Y(n2746) );
  CLKBUFX2TS U3270 ( .A(n67), .Y(n2771) );
  CLKBUFX2TS U3271 ( .A(n195), .Y(n2754) );
  INVXLTS U3272 ( .A(\addr_calc/N95 ), .Y(n195) );
  CLKBUFX2TS U3273 ( .A(n3), .Y(n2781) );
  CLKBUFX2TS U3274 ( .A(n259), .Y(n2745) );
  INVXLTS U3275 ( .A(\addr_calc/N63 ), .Y(n259) );
  CLKBUFX2TS U3276 ( .A(n67), .Y(n2773) );
  CLKBUFX2TS U3277 ( .A(n3), .Y(n2777) );
  CLKBUFX2TS U3278 ( .A(n323), .Y(n2737) );
  INVXLTS U3279 ( .A(\addr_calc/N9 ), .Y(n323) );
  CLKBUFX2TS U3280 ( .A(n67), .Y(n2769) );
  INVXLTS U3281 ( .A(\addr_calc/N159 ), .Y(n67) );
  CLKBUFX2TS U3282 ( .A(n3), .Y(n2779) );
  CLKBUFX2TS U3283 ( .A(n3), .Y(n2778) );
  INVXLTS U3284 ( .A(\addr_calc/N191 ), .Y(n3) );
  AO22X2TS U3285 ( .A0(n1822), .A1(\addr_calc/fir_read_calc/counter/N45 ), 
        .B0(n1673), .B1(n2004), .Y(n1096) );
  AO22X2TS U3286 ( .A0(n1151), .A1(\addr_calc/fir_read_calc/counter/N55 ), 
        .B0(n1674), .B1(n1994), .Y(n1086) );
  AO22X2TS U3287 ( .A0(n1824), .A1(\addr_calc/fir_read_calc/counter/N49 ), 
        .B0(n1671), .B1(n2001), .Y(n1092) );
  AO22X2TS U3288 ( .A0(n1827), .A1(\addr_calc/fir_read_calc/counter/N60 ), 
        .B0(n1671), .B1(n1884), .Y(n1081) );
  AO22X2TS U3289 ( .A0(n1823), .A1(\addr_calc/fir_read_calc/counter/N56 ), 
        .B0(n1674), .B1(n1893), .Y(n1085) );
  AO22X2TS U3290 ( .A0(n1824), .A1(\addr_calc/fir_read_calc/counter/N54 ), 
        .B0(n1743), .B1(n1895), .Y(n1087) );
  AO22X2TS U3291 ( .A0(n1825), .A1(\addr_calc/fir_read_calc/counter/N51 ), 
        .B0(n1673), .B1(n1997), .Y(n1090) );
  AO22X2TS U3292 ( .A0(n1827), .A1(\addr_calc/fir_read_calc/counter/N67 ), 
        .B0(n1663), .B1(\addr_calc/fir_read_calc/count[24] ), .Y(n1074) );
  AO22X2TS U3293 ( .A0(n1764), .A1(\addr_calc/fir_write_calc/counter/N46 ), 
        .B0(n1263), .B1(n1866), .Y(n1127) );
  AO22X2TS U3294 ( .A0(n1760), .A1(\addr_calc/fir_write_calc/counter/N51 ), 
        .B0(n1265), .B1(n1996), .Y(n1122) );
  AO22X2TS U3295 ( .A0(n1761), .A1(\addr_calc/fir_write_calc/counter/N54 ), 
        .B0(n1265), .B1(n1877), .Y(n1119) );
  AO22X2TS U3296 ( .A0(n1759), .A1(\addr_calc/fir_write_calc/counter/N48 ), 
        .B0(n1266), .B1(n1867), .Y(n1125) );
  AO22X2TS U3297 ( .A0(n1759), .A1(\addr_calc/fir_write_calc/counter/N49 ), 
        .B0(n1270), .B1(n1993), .Y(n1124) );
  AO22X2TS U3298 ( .A0(n1763), .A1(\addr_calc/fir_write_calc/counter/N56 ), 
        .B0(n1268), .B1(n1880), .Y(n1117) );
  AO22X2TS U3299 ( .A0(n1152), .A1(\addr_calc/fir_write_calc/counter/N70 ), 
        .B0(n1267), .B1(\addr_calc/fir_write_calc/count[27] ), .Y(n1103) );
  AO22X2TS U3300 ( .A0(n1760), .A1(\addr_calc/fir_write_calc/counter/N66 ), 
        .B0(n1259), .B1(n2563), .Y(n1107) );
  AO22X2TS U3301 ( .A0(n1763), .A1(\addr_calc/fir_write_calc/counter/N71 ), 
        .B0(n1262), .B1(n1896), .Y(n1102) );
  AO22X2TS U3302 ( .A0(n1760), .A1(\addr_calc/fir_write_calc/counter/N74 ), 
        .B0(n1262), .B1(n2550), .Y(n1099) );
  AO22X2TS U3303 ( .A0(n1752), .A1(\addr_calc/fft_read_calc/counter/N44 ), 
        .B0(n1979), .B1(n1475), .Y(n1033) );
  AO22X2TS U3304 ( .A0(n1754), .A1(\addr_calc/fft_read_calc/counter/N45 ), 
        .B0(n2056), .B1(n1477), .Y(n1032) );
  AO22X2TS U3305 ( .A0(n1761), .A1(\addr_calc/fir_write_calc/counter/N59 ), 
        .B0(n1264), .B1(n2564), .Y(n1114) );
  AO22X2TS U3306 ( .A0(n1759), .A1(\addr_calc/fir_write_calc/counter/N67 ), 
        .B0(n1264), .B1(n2577), .Y(n1106) );
  AO22X2TS U3307 ( .A0(n1152), .A1(\addr_calc/fir_write_calc/counter/N60 ), 
        .B0(\addr_calc/fir_write_calc/count[17] ), .B1(n1261), .Y(n1113) );
  AO22X2TS U3308 ( .A0(n1749), .A1(\addr_calc/fft_read_calc/counter/N46 ), 
        .B0(n2655), .B1(n1978), .Y(n1031) );
  AO22X2TS U3309 ( .A0(n1754), .A1(\addr_calc/fft_read_calc/counter/N51 ), 
        .B0(n2656), .B1(n2049), .Y(n1026) );
  AO22X2TS U3310 ( .A0(n1750), .A1(\addr_calc/fft_read_calc/counter/N52 ), 
        .B0(n2656), .B1(n2560), .Y(n1025) );
  AO22X2TS U3311 ( .A0(n1751), .A1(\addr_calc/fft_read_calc/counter/N53 ), 
        .B0(n2655), .B1(n1972), .Y(n1024) );
  AO22X2TS U3312 ( .A0(n1748), .A1(\addr_calc/fft_read_calc/counter/N48 ), 
        .B0(n2656), .B1(n1977), .Y(n1029) );
  AO22X2TS U3313 ( .A0(n1748), .A1(\addr_calc/fft_read_calc/counter/N68 ), 
        .B0(\addr_calc/fft_read_calc/count[25] ), .B1(n2659), .Y(n1009) );
  AO22X2TS U3314 ( .A0(n1752), .A1(\addr_calc/fft_read_calc/counter/N70 ), 
        .B0(\addr_calc/fft_read_calc/count[27] ), .B1(n2661), .Y(n1007) );
  AO22X2TS U3315 ( .A0(n1749), .A1(\addr_calc/fft_read_calc/counter/N66 ), 
        .B0(n2660), .B1(\addr_calc/fft_read_calc/count[23] ), .Y(n1011) );
  AO22X2TS U3316 ( .A0(n1750), .A1(\addr_calc/fft_read_calc/counter/N67 ), 
        .B0(n2658), .B1(\addr_calc/fft_read_calc/count[24] ), .Y(n1010) );
  AO22X2TS U3317 ( .A0(n1726), .A1(\addr_calc/fft_write_calc/counter/N68 ), 
        .B0(n2668), .B1(\addr_calc/fft_write_calc/count[25] ), .Y(n1041) );
  AO22X2TS U3318 ( .A0(n1753), .A1(\addr_calc/fft_read_calc/counter/N62 ), 
        .B0(n1956), .B1(n1477), .Y(n1015) );
  AO22X2TS U3319 ( .A0(n1722), .A1(\addr_calc/fft_write_calc/counter/N74 ), 
        .B0(n2662), .B1(\addr_calc/fft_write_calc/count[31] ), .Y(n1067) );
  AO22X2TS U3320 ( .A0(n1709), .A1(\addr_calc/iir_read_calc/counter/N45 ), 
        .B0(n2015), .B1(n2647), .Y(n969) );
  AO22X2TS U3321 ( .A0(n1714), .A1(\addr_calc/iir_read_calc/counter/N44 ), 
        .B0(n1898), .B1(n2647), .Y(n970) );
  AO22X2TS U3322 ( .A0(n1709), .A1(\addr_calc/iir_read_calc/counter/N71 ), 
        .B0(n2653), .B1(n2561), .Y(n943) );
  AO22X2TS U3323 ( .A0(n1710), .A1(\addr_calc/iir_read_calc/counter/N68 ), 
        .B0(n2650), .B1(\addr_calc/iir_read_calc/count[25] ), .Y(n946) );
  AO22X2TS U3324 ( .A0(n1713), .A1(\addr_calc/iir_read_calc/counter/N67 ), 
        .B0(\addr_calc/iir_read_calc/count[24] ), .B1(n2652), .Y(n947) );
  AO22X2TS U3325 ( .A0(n1709), .A1(\addr_calc/iir_read_calc/counter/N72 ), 
        .B0(n2653), .B1(n1840), .Y(n942) );
  AO22X2TS U3326 ( .A0(n1707), .A1(\addr_calc/iir_read_calc/counter/N59 ), 
        .B0(\addr_calc/iir_read_calc/count[16] ), .B1(n2647), .Y(n955) );
  AO22X2TS U3327 ( .A0(n1768), .A1(\addr_calc/iir_write_calc/counter/N47 ), 
        .B0(n2678), .B1(n1935), .Y(n998) );
  AO22X2TS U3328 ( .A0(n1769), .A1(\addr_calc/iir_write_calc/counter/N69 ), 
        .B0(n2678), .B1(n2573), .Y(n976) );
  AO22X2TS U3329 ( .A0(n1772), .A1(\addr_calc/iir_write_calc/counter/N70 ), 
        .B0(n2678), .B1(n1688), .Y(n975) );
  AO22X2TS U3330 ( .A0(n1770), .A1(\addr_calc/iir_write_calc/counter/N68 ), 
        .B0(n2678), .B1(\addr_calc/iir_write_calc/count[25] ), .Y(n977) );
  AO22X2TS U3331 ( .A0(n1769), .A1(\addr_calc/iir_write_calc/counter/N73 ), 
        .B0(n2672), .B1(n1854), .Y(n1003) );
  AO22X2TS U3332 ( .A0(n1770), .A1(\addr_calc/iir_write_calc/counter/N62 ), 
        .B0(n2672), .B1(\addr_calc/iir_write_calc/count[19] ), .Y(n983) );
  CLKBUFX2TS U3333 ( .A(data_from_iir), .Y(n2718) );
  CLKBUFX2TS U3334 ( .A(n451), .Y(n2721) );
  CLKBUFX2TS U3335 ( .A(n451), .Y(n2722) );
  CLKBUFX2TS U3336 ( .A(n451), .Y(n2723) );
  CLKBUFX2TS U3337 ( .A(n2645), .Y(n2750) );
  CLKBUFX2TS U3338 ( .A(n2644), .Y(n2758) );
  CLKBUFX2TS U3339 ( .A(n2643), .Y(n2766) );
  CLKBUFX2TS U3340 ( .A(n2641), .Y(n2782) );
  CLKBUFX2TS U3341 ( .A(data_from_iir), .Y(n2717) );
  CLKBUFX2TS U3342 ( .A(n2646), .Y(n2740) );
  CLKBUFX2TS U3343 ( .A(n2646), .Y(n2742) );
  CLKBUFX2TS U3344 ( .A(n2645), .Y(n2748) );
  CLKBUFX2TS U3345 ( .A(n2644), .Y(n2756) );
  CLKBUFX2TS U3346 ( .A(data_to_fir), .Y(n2708) );
  CLKBUFX2TS U3347 ( .A(n515), .Y(n2709) );
  CLKBUFX2TS U3348 ( .A(n515), .Y(n2712) );
  CLKBUFX2TS U3349 ( .A(n515), .Y(n2713) );
  CLKBUFX2TS U3350 ( .A(data_to_iir), .Y(n2726) );
  CLKBUFX2TS U3351 ( .A(n387), .Y(n2727) );
  CLKBUFX2TS U3352 ( .A(data_to_fft), .Y(n2690) );
  CLKBUFX2TS U3353 ( .A(n387), .Y(n2730) );
  CLKBUFX2TS U3354 ( .A(n387), .Y(n2731) );
  CLKBUFX2TS U3355 ( .A(data_from_fft), .Y(n2681) );
  CLKBUFX2TS U3356 ( .A(data_from_fft), .Y(n2682) );
  CLKBUFX2TS U3357 ( .A(n707), .Y(n2685) );
  CLKBUFX2TS U3358 ( .A(n707), .Y(n2686) );
  CLKBUFX2TS U3359 ( .A(n707), .Y(n2687) );
  CLKBUFX2TS U3360 ( .A(data_from_fir), .Y(n2699) );
  CLKBUFX2TS U3361 ( .A(data_from_fir), .Y(n2700) );
  CLKBUFX2TS U3362 ( .A(n579), .Y(n2703) );
  CLKBUFX2TS U3363 ( .A(n579), .Y(n2704) );
  CLKBUFX2TS U3364 ( .A(n579), .Y(n2705) );
  CLKBUFX2TS U3365 ( .A(n2643), .Y(n2764) );
  CLKBUFX2TS U3366 ( .A(n2643), .Y(n2759) );
  CLKBUFX2TS U3367 ( .A(n2641), .Y(n2775) );
  CLKBUFX2TS U3368 ( .A(n2645), .Y(n2743) );
  CLKBUFX2TS U3369 ( .A(n2646), .Y(n2735) );
  CLKBUFX2TS U3370 ( .A(n2642), .Y(n2772) );
  CLKBUFX2TS U3371 ( .A(n2641), .Y(n2780) );
  CLKBUFX2TS U3372 ( .A(n2646), .Y(n2736) );
  CLKBUFX2TS U3373 ( .A(n2642), .Y(n2767) );
  CLKBUFX2TS U3374 ( .A(n2645), .Y(n2744) );
  CLKBUFX2TS U3375 ( .A(n2642), .Y(n2768) );
  CLKBUFX2TS U3376 ( .A(n2642), .Y(n2774) );
  CLKBUFX2TS U3377 ( .A(n2643), .Y(n2760) );
  CLKBUFX2TS U3378 ( .A(n2641), .Y(n2776) );
  CLKBUFX2TS U3379 ( .A(n2644), .Y(n2752) );
  CLKBUFX2TS U3380 ( .A(n2644), .Y(n2751) );
  CLKBUFX2TS U3381 ( .A(n643), .Y(n2691) );
  CLKBUFX2TS U3382 ( .A(n643), .Y(n2694) );
  CLKBUFX2TS U3383 ( .A(n643), .Y(n2695) );
  OAI21XLTS U3384 ( .A0(n2810), .A1(n2808), .B0(fir_enable), .Y(n2811) );
  OAI21XLTS U3385 ( .A0(\addr_calc/fir_write_calc/counter/N43 ), .A1(n2804), 
        .B0(n2069), .Y(n2806) );
  NAND4X1TS U3386 ( .A(n880), .B(n881), .C(n882), .D(n883), .Y(n2800) );
  NAND4X1TS U3387 ( .A(n861), .B(n862), .C(n863), .D(n864), .Y(n2801) );
  NOR4XLTS U3388 ( .A(n1872), .B(n1995), .C(
        \addr_calc/fir_write_calc/count[7] ), .D(n1992), .Y(n862) );
  NAND4X1TS U3389 ( .A(n865), .B(n866), .C(n867), .D(n868), .Y(n2802) );
  NOR4XLTS U3390 ( .A(n2560), .B(n2049), .C(\addr_calc/fft_read_calc/count[7] ), .D(n2052), .Y(n829) );
  NOR4XLTS U3391 ( .A(n1936), .B(n2026), .C(n1934), .D(n2030), .Y(n843) );
  NAND4X1TS U3392 ( .A(n810), .B(n811), .C(n812), .D(n813), .Y(n2783) );
  NOR4XLTS U3393 ( .A(\addr_calc/iir_read_calc/count[9] ), .B(n2583), .C(
        \addr_calc/iir_read_calc/count[7] ), .D(n2018), .Y(n811) );
  NAND4X1TS U3394 ( .A(n814), .B(n815), .C(n816), .D(n817), .Y(n2784) );
  NAND4X1TS U3395 ( .A(n915), .B(n916), .C(n917), .D(n918), .Y(n2788) );
  NOR4XLTS U3396 ( .A(n2562), .B(n2041), .C(
        \addr_calc/iir_write_calc/count[7] ), .D(n2039), .Y(n916) );
  NAND4X1TS U3397 ( .A(n919), .B(n920), .C(n921), .D(n922), .Y(n2789) );
endmodule

