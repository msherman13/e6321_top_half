library verilog;
use verilog.vl_types.all;
entity TIEHITS is
    port(
        Y               : out    vl_logic
    );
end TIEHITS;
