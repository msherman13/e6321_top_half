library verilog;
use verilog.vl_types.all;
entity DLY2X4TS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end DLY2X4TS;
