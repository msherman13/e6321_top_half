

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO top_level 
  PIN acc_fft_data_out[31] 
  END acc_fft_data_out[31]
  PIN acc_fft_data_out[30] 
  END acc_fft_data_out[30]
  PIN acc_fft_data_out[29] 
  END acc_fft_data_out[29]
  PIN acc_fft_data_out[28] 
  END acc_fft_data_out[28]
  PIN acc_fft_data_out[27] 
  END acc_fft_data_out[27]
  PIN acc_fft_data_out[26] 
  END acc_fft_data_out[26]
  PIN acc_fft_data_out[25] 
  END acc_fft_data_out[25]
  PIN acc_fft_data_out[24] 
  END acc_fft_data_out[24]
  PIN acc_fft_data_out[23] 
  END acc_fft_data_out[23]
  PIN acc_fft_data_out[22] 
  END acc_fft_data_out[22]
  PIN acc_fft_data_out[21] 
  END acc_fft_data_out[21]
  PIN acc_fft_data_out[20] 
  END acc_fft_data_out[20]
  PIN acc_fft_data_out[19] 
  END acc_fft_data_out[19]
  PIN acc_fft_data_out[18] 
  END acc_fft_data_out[18]
  PIN acc_fft_data_out[17] 
  END acc_fft_data_out[17]
  PIN acc_fft_data_out[16] 
  END acc_fft_data_out[16]
  PIN acc_fft_data_out[15] 
  END acc_fft_data_out[15]
  PIN acc_fft_data_out[14] 
  END acc_fft_data_out[14]
  PIN acc_fft_data_out[13] 
  END acc_fft_data_out[13]
  PIN acc_fft_data_out[12] 
  END acc_fft_data_out[12]
  PIN acc_fft_data_out[11] 
  END acc_fft_data_out[11]
  PIN acc_fft_data_out[10] 
  END acc_fft_data_out[10]
  PIN acc_fft_data_out[9] 
  END acc_fft_data_out[9]
  PIN acc_fft_data_out[8] 
  END acc_fft_data_out[8]
  PIN acc_fft_data_out[7] 
  END acc_fft_data_out[7]
  PIN acc_fft_data_out[6] 
  END acc_fft_data_out[6]
  PIN acc_fft_data_out[5] 
  END acc_fft_data_out[5]
  PIN acc_fft_data_out[4] 
  END acc_fft_data_out[4]
  PIN acc_fft_data_out[3] 
  END acc_fft_data_out[3]
  PIN acc_fft_data_out[2] 
  END acc_fft_data_out[2]
  PIN acc_fft_data_out[1] 
  END acc_fft_data_out[1]
  PIN acc_fft_data_out[0] 
  END acc_fft_data_out[0]
  PIN acc_fft_data_in[31] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 36.0045 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[31]
  PIN acc_fft_data_in[30] 
    ANTENNAPARTIALMETALAREA 3.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 37.8063 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 140.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[30]
  PIN acc_fft_data_in[29] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 21.1396 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 75.5225 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.95495 LAYER VQ ;
  END acc_fft_data_in[29]
  PIN acc_fft_data_in[28] 
    ANTENNAPARTIALMETALAREA 3.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.3108 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 157.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[28]
  PIN acc_fft_data_in[27] 
    ANTENNAPARTIALMETALAREA 3.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 37.8063 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 140.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[27]
  PIN acc_fft_data_in[26] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[26]
  PIN acc_fft_data_in[25] 
    ANTENNAPARTIALMETALAREA 43.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 159.914 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.7162 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END acc_fft_data_in[25]
  PIN acc_fft_data_in[24] 
    ANTENNAPARTIALMETALAREA 5.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.978 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.0225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END acc_fft_data_in[24]
  PIN acc_fft_data_in[23] 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 27.8964 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 103.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[23]
  PIN acc_fft_data_in[22] 
    ANTENNAPARTIALMETALAREA 3.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.3108 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 157.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[22]
  PIN acc_fft_data_in[21] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[21]
  PIN acc_fft_data_in[20] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[20]
  PIN acc_fft_data_in[19] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 54.9234 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 208.856 LAYER MQ ;
    ANTENNAMAXCUTCAR 3.15315 LAYER VQ ;
  END acc_fft_data_in[19]
  PIN acc_fft_data_in[18] 
    ANTENNAPARTIALMETALAREA 3.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.3108 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 157.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[18]
  PIN acc_fft_data_in[17] 
    ANTENNAPARTIALMETALAREA 12.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 46.25 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.3829 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 149.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fft_data_in[17]
  PIN acc_fft_data_in[16] 
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 119.563 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 446.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fft_data_in[16]
  PIN acc_fft_data_in[15] 
    ANTENNAPARTIALMETALAREA 3.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 39.6081 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 147.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[15]
  PIN acc_fft_data_in[14] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[14]
  PIN acc_fft_data_in[13] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[13]
  PIN acc_fft_data_in[12] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[12]
  PIN acc_fft_data_in[11] 
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 58.527 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 217.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[11]
  PIN acc_fft_data_in[10] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 36.0045 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[10]
  PIN acc_fft_data_in[9] 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 27.8964 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 103.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[9]
  PIN acc_fft_data_in[8] 
    ANTENNAPARTIALMETALAREA 4.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.834 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 55.3739 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 207.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[8]
  PIN acc_fft_data_in[7] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 74.2928 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 285.523 LAYER MQ ;
    ANTENNAMAXCUTCAR 3.15315 LAYER VQ ;
  END acc_fft_data_in[7]
  PIN acc_fft_data_in[6] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 36.0045 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[6]
  PIN acc_fft_data_in[5] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 31.5 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 112.189 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.95495 LAYER VQ ;
  END acc_fft_data_in[5]
  PIN acc_fft_data_in[4] 
    ANTENNAPARTIALMETALAREA 1.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.514 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 92.648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2136 LAYER M3 ; 
    ANTENNAMAXAREACAR 116.96 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 438.586 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.561798 LAYER VL ;
  END acc_fft_data_in[4]
  PIN acc_fft_data_in[3] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[3]
  PIN acc_fft_data_in[2] 
    ANTENNAPARTIALMETALAREA 15.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 55.722 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.136 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.3829 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 156.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fft_data_in[2]
  PIN acc_fft_data_in[1] 
    ANTENNAPARTIALMETALAREA 4.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.65 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 52.2207 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 193.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fft_data_in[1]
  PIN acc_fft_data_in[0] 
    ANTENNAPARTIALMETALAREA 3.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.8604 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fft_data_in[0]
  PIN acc_fir_data_out[31] 
  END acc_fir_data_out[31]
  PIN acc_fir_data_out[30] 
  END acc_fir_data_out[30]
  PIN acc_fir_data_out[29] 
  END acc_fir_data_out[29]
  PIN acc_fir_data_out[28] 
  END acc_fir_data_out[28]
  PIN acc_fir_data_out[27] 
  END acc_fir_data_out[27]
  PIN acc_fir_data_out[26] 
  END acc_fir_data_out[26]
  PIN acc_fir_data_out[25] 
  END acc_fir_data_out[25]
  PIN acc_fir_data_out[24] 
  END acc_fir_data_out[24]
  PIN acc_fir_data_out[23] 
  END acc_fir_data_out[23]
  PIN acc_fir_data_out[22] 
  END acc_fir_data_out[22]
  PIN acc_fir_data_out[21] 
  END acc_fir_data_out[21]
  PIN acc_fir_data_out[20] 
  END acc_fir_data_out[20]
  PIN acc_fir_data_out[19] 
  END acc_fir_data_out[19]
  PIN acc_fir_data_out[18] 
  END acc_fir_data_out[18]
  PIN acc_fir_data_out[17] 
  END acc_fir_data_out[17]
  PIN acc_fir_data_out[16] 
  END acc_fir_data_out[16]
  PIN acc_fir_data_out[15] 
  END acc_fir_data_out[15]
  PIN acc_fir_data_out[14] 
  END acc_fir_data_out[14]
  PIN acc_fir_data_out[13] 
  END acc_fir_data_out[13]
  PIN acc_fir_data_out[12] 
  END acc_fir_data_out[12]
  PIN acc_fir_data_out[11] 
  END acc_fir_data_out[11]
  PIN acc_fir_data_out[10] 
  END acc_fir_data_out[10]
  PIN acc_fir_data_out[9] 
  END acc_fir_data_out[9]
  PIN acc_fir_data_out[8] 
  END acc_fir_data_out[8]
  PIN acc_fir_data_out[7] 
  END acc_fir_data_out[7]
  PIN acc_fir_data_out[6] 
  END acc_fir_data_out[6]
  PIN acc_fir_data_out[5] 
  END acc_fir_data_out[5]
  PIN acc_fir_data_out[4] 
  END acc_fir_data_out[4]
  PIN acc_fir_data_out[3] 
  END acc_fir_data_out[3]
  PIN acc_fir_data_out[2] 
  END acc_fir_data_out[2]
  PIN acc_fir_data_out[1] 
  END acc_fir_data_out[1]
  PIN acc_fir_data_out[0] 
  END acc_fir_data_out[0]
  PIN acc_fir_data_in[31] 
    ANTENNAPARTIALMETALAREA 27.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 100.714 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.8604 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[31]
  PIN acc_fir_data_in[30] 
    ANTENNAPARTIALMETALAREA 2.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 108.302 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 409.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[30]
  PIN acc_fir_data_in[29] 
    ANTENNAPARTIALMETALAREA 1.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.586 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.352 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 65.0586 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 246.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[29]
  PIN acc_fir_data_in[28] 
    ANTENNAPARTIALMETALAREA 6.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 98.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 373.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[28]
  PIN acc_fir_data_in[27] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 155.824 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 582.189 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.7027 LAYER VQ ;
  END acc_fir_data_in[27]
  PIN acc_fir_data_in[26] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 47.7162 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 175.523 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.95495 LAYER VQ ;
  END acc_fir_data_in[26]
  PIN acc_fir_data_in[25] 
    ANTENNAPARTIALMETALAREA 5.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.018 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.04 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 107.851 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 409.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[25]
  PIN acc_fir_data_in[24] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.0856 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 163.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[24]
  PIN acc_fir_data_in[23] 
    ANTENNAPARTIALMETALAREA 3.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.3108 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 157.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[23]
  PIN acc_fir_data_in[22] 
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 58.527 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 217.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[22]
  PIN acc_fir_data_in[21] 
    ANTENNAPARTIALMETALAREA 5.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.314 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 60.3288 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 223.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[21]
  PIN acc_fir_data_in[20] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 36.0045 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[20]
  PIN acc_fir_data_in[19] 
    ANTENNAPARTIALMETALAREA 19.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 73.778 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.24775 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 19.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END acc_fir_data_in[19]
  PIN acc_fir_data_in[18] 
    ANTENNAPARTIALMETALAREA 3.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 37.8063 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 140.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[18]
  PIN acc_fir_data_in[17] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[17]
  PIN acc_fir_data_in[16] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[16]
  PIN acc_fir_data_in[15] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 42.3108 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 152.189 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.95495 LAYER VQ ;
  END acc_fir_data_in[15]
  PIN acc_fir_data_in[14] 
    ANTENNAPARTIALMETALAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.642 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 76.545 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 283.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[14]
  PIN acc_fir_data_in[13] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[13]
  PIN acc_fir_data_in[12] 
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 58.527 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 217.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[12]
  PIN acc_fir_data_in[11] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[11]
  PIN acc_fir_data_in[10] 
    ANTENNAPARTIALMETALAREA 2.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.9955 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 100.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END acc_fir_data_in[10]
  PIN acc_fir_data_in[9] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 31.5 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 112.189 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.95495 LAYER VQ ;
  END acc_fir_data_in[9]
  PIN acc_fir_data_in[8] 
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.1577 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 56.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[8]
  PIN acc_fir_data_in[7] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 111.005 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 416.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[7]
  PIN acc_fir_data_in[6] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 96.5901 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 366.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[6]
  PIN acc_fir_data_in[5] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.1847 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 163.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END acc_fir_data_in[5]
  PIN acc_fir_data_in[4] 
    ANTENNAPARTIALMETALAREA 11.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 43.882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1056 LAYER M3 ; 
    ANTENNAMAXAREACAR 61.5417 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 231.644 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.51515 LAYER VL ;
  END acc_fir_data_in[4]
  PIN acc_fir_data_in[3] 
    ANTENNAPARTIALMETALAREA 12.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 46.546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 143.887 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 536.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[3]
  PIN acc_fir_data_in[2] 
    ANTENNAPARTIALMETALAREA 10.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 40.33 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 56.9505 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 219.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[2]
  PIN acc_fir_data_in[1] 
    ANTENNAPARTIALMETALAREA 13.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 51.578 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 47.0405 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 179.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[1]
  PIN acc_fir_data_in[0] 
    ANTENNAPARTIALMETALAREA 16.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.938 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 70.464 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 266.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_data_in[0]
  PIN addr[31] 
    ANTENNAPARTIALMETALAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.642 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 75.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.90451 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.7408 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL ;
  END addr[31]
  PIN addr[30] 
    ANTENNAPARTIALMETALAREA 1.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.106 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.76 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.38214 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.02438 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[30]
  PIN addr[29] 
    ANTENNAPARTIALMETALAREA 11.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 44.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.98029 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.24375 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL ;
  END addr[29]
  PIN addr[28] 
    ANTENNAPARTIALMETALAREA 15.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.906 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.52311 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.48796 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL ;
  END addr[28]
  PIN addr[27] 
    ANTENNAPARTIALMETALAREA 12.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 44.474 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.69711 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 13.4747 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.88 LAYER M3 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.28931 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.6872 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0617284 LAYER VL ;
  END addr[27]
  PIN addr[26] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER MQ ; 
    ANTENNAMAXAREACAR 3.96813 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 14.5488 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.108025 LAYER VQ ;
  END addr[26]
  PIN addr[25] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.40313 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.2083 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL ;
  END addr[25]
  PIN addr[24] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.64988 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.06605 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL ;
  END addr[24]
  PIN addr[23] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER MQ ; 
    ANTENNAMAXAREACAR 1.29244 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 4.77197 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.100309 LAYER VQ ;
  END addr[23]
  PIN addr[22] 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.922 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.72 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.42303 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.14514 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[22]
  PIN addr[21] 
    ANTENNAPARTIALMETALAREA 4.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.14309 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.07477 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0578704 LAYER VL ;
  END addr[21]
  PIN addr[20] 
    ANTENNAPARTIALMETALAREA 6.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.866 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.97257 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.22234 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER M3 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.37959 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.74973 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[20]
  PIN addr[19] 
    ANTENNAPARTIALMETALAREA 1.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.106 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.82967 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.68642 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[19]
  PIN addr[18] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.19248 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.02886 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[18]
  PIN addr[17] 
    ANTENNAPARTIALMETALAREA 4.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.466 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.00058 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.32994 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL ;
  END addr[17]
  PIN addr[16] 
    ANTENNAPARTIALMETALAREA 4.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.65 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.912 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.858565 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.01487 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 68.672 LAYER M3 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.74784 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.3266 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[16]
  PIN addr[15] 
    ANTENNAPARTIALMETALAREA 1.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.514 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.05035 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.5294 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[15]
  PIN addr[14] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER MQ ; 
    ANTENNAMAXAREACAR 2.26408 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 8.29271 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.100309 LAYER VQ ;
  END addr[14]
  PIN addr[13] 
    ANTENNAPARTIALMETALAREA 2.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.60613 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.87253 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL ;
  END addr[13]
  PIN addr[12] 
    ANTENNAPARTIALMETALAREA 5.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.202 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.78738 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.4515 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.352 LAYER M3 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.49919 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.12087 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[12]
  PIN addr[11] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER MQ ; 
    ANTENNAMAXAREACAR 3.00887 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 11.0586 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.123457 LAYER VQ ;
  END addr[11]
  PIN addr[10] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.27334 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.72577 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[10]
  PIN addr[9] 
    ANTENNAPARTIALMETALAREA 1.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.29 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.11262 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.4262 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[9]
  PIN addr[8] 
    ANTENNAPARTIALMETALAREA 1.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.994 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.61223 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.2677 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL ;
  END addr[8]
  PIN addr[7] 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 68.376 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.28669 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.39259 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL ;
  END addr[7]
  PIN addr[6] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.8684 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.78696 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.115741 LAYER VL ;
  END addr[6]
  PIN addr[5] 
    ANTENNAPARTIALMETALAREA 7.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.12 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.008 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.91107 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.00085 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[5]
  PIN addr[4] 
    ANTENNAPARTIALMETALAREA 0.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.33 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 68.968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.3532 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 12.5568 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VL ;
  END addr[4]
  PIN addr[3] 
    ANTENNAPARTIALMETALAREA 0.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.554 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 72.224 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.64834 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.95841 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL ;
  END addr[3]
  PIN addr[2] 
    ANTENNAPARTIALMETALAREA 11.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 42.106 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.28067 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.63164 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0578704 LAYER VL ;
  END addr[2]
  PIN addr[1] 
    ANTENNAPARTIALMETALAREA 8.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.338 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.136 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.81424 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.5865 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VL ;
  END addr[1]
  PIN addr[0] 
    ANTENNAPARTIALMETALAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 20.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.85783 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.75085 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0694444 LAYER VL ;
  END addr[0]
  PIN data_bus[31] 
    ANTENNAPARTIALMETALAREA 3.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.49363 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.1706 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[31]
  PIN data_bus[30] 
    ANTENNAPARTIALMETALAREA 4.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.948 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.29688 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.52824 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[30]
  PIN data_bus[29] 
    ANTENNAPARTIALMETALAREA 5.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.978 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.82002 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.70069 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[29]
  PIN data_bus[28] 
    ANTENNAPARTIALMETALAREA 10.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 37.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.20289 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.37454 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[28]
  PIN data_bus[27] 
    ANTENNAPARTIALMETALAREA 20.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 76.738 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.3397 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 23.3888 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[27]
  PIN data_bus[26] 
    ANTENNAPARTIALMETALAREA 17.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 63.418 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 5.17859 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 18.9561 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[26]
  PIN data_bus[25] 
    ANTENNAPARTIALMETALAREA 12.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 44.474 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.93762 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 14.469 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[25]
  PIN data_bus[24] 
    ANTENNAPARTIALMETALAREA 12.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 44.474 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.69271 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.23773 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[24]
  PIN data_bus[23] 
    ANTENNAPARTIALMETALAREA 4.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.762 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.45174 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.16678 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[23]
  PIN data_bus[22] 
    ANTENNAPARTIALMETALAREA 3.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.4022 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.06701 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[22]
  PIN data_bus[21] 
    ANTENNAPARTIALMETALAREA 3.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.2434 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 4.39595 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[21]
  PIN data_bus[20] 
    ANTENNAPARTIALMETALAREA 4.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.426 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.66007 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.93762 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[20]
  PIN data_bus[19] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.89641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 18.0711 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[19]
  PIN data_bus[18] 
    ANTENNAPARTIALMETALAREA 5.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.09 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.8684 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.70845 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[18]
  PIN data_bus[17] 
    ANTENNAPARTIALMETALAREA 6.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.37326 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.73542 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[17]
  PIN data_bus[16] 
    ANTENNAPARTIALMETALAREA 4.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.834 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.63808 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.68472 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[16]
  PIN data_bus[15] 
    ANTENNAPARTIALMETALAREA 2.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.434 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.03507 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.62512 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[15]
  PIN data_bus[14] 
    ANTENNAPARTIALMETALAREA 4.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.762 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.45174 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.16678 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[14]
  PIN data_bus[13] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.826736 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.85428 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[13]
  PIN data_bus[12] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ ; 
    ANTENNAMAXAREACAR 0.629977 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 2.04063 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VQ ;
  END data_bus[12]
  PIN data_bus[11] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.826736 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.85428 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[11]
  PIN data_bus[10] 
    ANTENNAPARTIALMETALAREA 4.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.058 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.52488 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.43738 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[10]
  PIN data_bus[9] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.826736 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.85428 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0231481 LAYER V2 ;
  END data_bus[9]
  PIN data_bus[8] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ ; 
    ANTENNAMAXAREACAR 1.19711 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 4.09618 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VQ ;
  END data_bus[8]
  PIN data_bus[7] 
    ANTENNAPARTIALMETALAREA 2.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.73 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.07234 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.0016 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[7]
  PIN data_bus[6] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ ; 
    ANTENNAMAXAREACAR 1.00174 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 3.66076 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VQ ;
  END data_bus[6]
  PIN data_bus[5] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ ; 
    ANTENNAMAXAREACAR 2.23877 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 8.20729 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VQ ;
  END data_bus[5]
  PIN data_bus[4] 
    ANTENNAPARTIALMETALAREA 4.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.43438 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.31667 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[4]
  PIN data_bus[3] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.17419 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.97847 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[3]
  PIN data_bus[2] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ ; 
    ANTENNAMAXAREACAR 3.211 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 11.6332 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VQ ;
  END data_bus[2]
  PIN data_bus[1] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER MQ ; 
    ANTENNAMAXAREACAR 6.19711 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 22.5962 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.138889 LAYER VQ ;
  END data_bus[1]
  PIN data_bus[0] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.456 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.03854 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 14.8236 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0462963 LAYER VL ;
  END data_bus[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.576 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7016 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.89563 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.3162 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0470146 LAYER VL ;
  END clk
  PIN reset 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 50.4189 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 185.523 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.95495 LAYER VQ ;
  END reset
  PIN acc_fft_get 
    ANTENNAPARTIALMETALAREA 8.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.042 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.7342 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 156.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fft_get
  PIN acc_fft_put 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 65.2838 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 248.856 LAYER MQ ;
    ANTENNAMAXCUTCAR 3.15315 LAYER VQ ;
  END acc_fft_put
  PIN acc_fir_get 
    ANTENNAPARTIALMETALAREA 3.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_get
  PIN acc_fir_put 
    ANTENNAPARTIALMETALAREA 5.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.682 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 114.608 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 436.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END acc_fir_put
  PIN fft_enable 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7272 LAYER MQ ; 
    ANTENNAMAXAREACAR 23.6574 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 88.4455 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.892307 LAYER VQ ;
  END fft_enable
  PIN fir_enable 
    ANTENNAPARTIALMETALAREA 19.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 71.706 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M2 ; 
    ANTENNAMAXAREACAR 133.833 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 496.976 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.728 LAYER M3 ;
    ANTENNAGATEAREA 4.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 137.06 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 509.06 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END fir_enable
  PIN to_fft_empty 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.16 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.5808 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.8147 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 52.3224 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.806452 LAYER VL ;
  END to_fft_empty
  PIN from_fft_full 
    ANTENNAPARTIALMETALAREA 11.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 42.994 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.62364 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.56523 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER VL ;
  END from_fft_full
  PIN to_fir_empty 
    ANTENNAPARTIALMETALAREA 7.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.01 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.5328 LAYER M3 ; 
    ANTENNAMAXAREACAR 92.242 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 340.974 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.98413 LAYER VL ;
  END to_fir_empty
  PIN from_fir_full 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER MQ ; 
    ANTENNAMAXAREACAR 4.68432 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 17.0706 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.136364 LAYER VQ ;
  END from_fir_full
  PIN ram_read_enable 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.207 LAYER MQ ; 
    ANTENNAMAXAREACAR 1.55162 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 5.29591 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0666019 LAYER VQ ;
  END ram_read_enable
  PIN ram_write_enable 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.898 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.938854 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.46253 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0138026 LAYER V2 ;
  END ram_write_enable
END top_level

END LIBRARY
