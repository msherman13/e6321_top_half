library verilog;
use verilog.vl_types.all;
entity BUFX2TS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end BUFX2TS;
