module top_level (
	clk, 
	reset, 
	acc_fft_get, 
	acc_fft_put, 
	acc_fir_get, 
	acc_fir_put, 
	acc_fft_data_out, 
	acc_fft_data_in, 
	acc_fir_data_out, 
	acc_fir_data_in, 
	fft_enable, 
	fir_enable, 
	to_fft_empty, 
	from_fft_full, 
	to_fir_empty, 
	from_fir_full, 
	ram_read_enable, 
	ram_write_enable, 
	addr, 
	data_bus);
   input clk;
   input reset;
   input acc_fft_get;
   input acc_fft_put;
   input acc_fir_get;
   input acc_fir_put;
   input [31:0] acc_fft_data_out;
   input [31:0] acc_fft_data_in;
   input [31:0] acc_fir_data_out;
   input [31:0] acc_fir_data_in;
   output fft_enable;
   output fir_enable;
   output to_fft_empty;
   output from_fft_full;
   output to_fir_empty;
   output from_fir_full;
   output ram_read_enable;
   output ram_write_enable;
   output [31:0] addr;
   inout [31:0] data_bus;

   // Internal wires
   wire clk__L1_N0;
   wire FE_OFN1825_n7107;
   wire FE_OFN1824_router_addr_calc_fir_read_calc_count_5_;
   wire FE_OFN1823_n4643;
   wire FE_OFN1822_n4643;
   wire FE_OFN1821_acc_fft_data_in_28_;
   wire FE_OFN1820_acc_fft_data_in_28_;
   wire FE_OFN1819_acc_fft_data_in_28_;
   wire FE_OFN1818_acc_fir_data_in_26_;
   wire FE_MDBN15_;
   wire FE_OFN1817_acc_fir_data_in_0_;
   wire FE_OFN1816_acc_fir_data_in_0_;
   wire FE_OFN1815_acc_fir_data_in_0_;
   wire FE_OFN1814_acc_fir_data_in_0_;
   wire FE_OFN1813_acc_fir_data_in_0_;
   wire FE_OFN1812_acc_fir_data_in_0_;
   wire FE_OFN1811_acc_fir_data_in_0_;
   wire FE_OFN1810_acc_fir_data_in_0_;
   wire FE_OFN1809_acc_fir_data_in_0_;
   wire FE_OFN1808_acc_fir_data_in_0_;
   wire FE_OFN1807_acc_fir_data_in_1_;
   wire FE_OFN1806_acc_fir_data_in_1_;
   wire FE_OFN1805_acc_fir_data_in_1_;
   wire FE_OFN1804_acc_fir_data_in_1_;
   wire FE_OFN1803_acc_fir_data_in_1_;
   wire FE_OFN1802_acc_fir_data_in_1_;
   wire FE_OFN1801_acc_fir_data_in_2_;
   wire FE_OFN1800_acc_fir_data_in_2_;
   wire FE_OFN1799_acc_fir_data_in_2_;
   wire FE_OFN1798_acc_fir_data_in_2_;
   wire FE_OFN1797_acc_fir_data_in_2_;
   wire FE_OFN1796_acc_fir_data_in_2_;
   wire FE_OFN1795_acc_fir_data_in_2_;
   wire FE_OFN1794_acc_fir_data_in_3_;
   wire FE_OFN1793_acc_fir_data_in_3_;
   wire FE_OFN1792_acc_fir_data_in_3_;
   wire FE_OFN1791_acc_fir_data_in_3_;
   wire FE_OFN1790_acc_fir_data_in_3_;
   wire FE_OFN1789_acc_fir_data_in_4_;
   wire FE_OFN1788_acc_fir_data_in_4_;
   wire FE_OFN1787_acc_fir_data_in_4_;
   wire FE_OFN1786_acc_fir_data_in_4_;
   wire FE_OFN1785_acc_fir_data_in_4_;
   wire FE_OFN1784_acc_fir_data_in_4_;
   wire FE_OFN1783_acc_fir_data_in_4_;
   wire FE_OFN1782_acc_fir_data_in_5_;
   wire FE_OFN1781_acc_fir_data_in_5_;
   wire FE_OFN1780_acc_fir_data_in_5_;
   wire FE_OFN1779_acc_fir_data_in_5_;
   wire FE_OFN1778_acc_fir_data_in_5_;
   wire FE_OFN1777_acc_fir_data_in_5_;
   wire FE_OFN1776_acc_fir_data_in_6_;
   wire FE_OFN1775_acc_fir_data_in_6_;
   wire FE_OFN1774_acc_fir_data_in_6_;
   wire FE_OFN1773_acc_fir_data_in_6_;
   wire FE_OFN1772_acc_fir_data_in_6_;
   wire FE_OFN1771_acc_fir_data_in_6_;
   wire FE_OFN1770_acc_fir_data_in_6_;
   wire FE_OFN1769_acc_fir_data_in_6_;
   wire FE_OFN1768_acc_fir_data_in_7_;
   wire FE_OFN1767_acc_fir_data_in_7_;
   wire FE_OFN1766_acc_fir_data_in_7_;
   wire FE_OFN1765_acc_fir_data_in_7_;
   wire FE_OFN1764_acc_fir_data_in_7_;
   wire FE_OFN1763_acc_fir_data_in_7_;
   wire FE_OFN1762_acc_fir_data_in_7_;
   wire FE_OFN1761_acc_fir_data_in_8_;
   wire FE_OFN1760_acc_fir_data_in_8_;
   wire FE_OFN1759_acc_fir_data_in_8_;
   wire FE_OFN1758_acc_fir_data_in_8_;
   wire FE_OFN1757_acc_fir_data_in_8_;
   wire FE_OFN1756_acc_fir_data_in_8_;
   wire FE_OFN1755_acc_fir_data_in_9_;
   wire FE_OFN1754_acc_fir_data_in_9_;
   wire FE_OFN1753_acc_fir_data_in_9_;
   wire FE_OFN1752_acc_fir_data_in_9_;
   wire FE_OFN1751_acc_fir_data_in_9_;
   wire FE_OFN1750_acc_fir_data_in_10_;
   wire FE_OFN1749_acc_fir_data_in_10_;
   wire FE_OFN1748_acc_fir_data_in_10_;
   wire FE_OFN1747_acc_fir_data_in_10_;
   wire FE_OFN1746_acc_fir_data_in_10_;
   wire FE_OFN1745_acc_fir_data_in_11_;
   wire FE_OFN1744_acc_fir_data_in_11_;
   wire FE_OFN1743_acc_fir_data_in_11_;
   wire FE_OFN1742_acc_fir_data_in_11_;
   wire FE_OFN1741_acc_fir_data_in_11_;
   wire FE_OFN1740_acc_fir_data_in_12_;
   wire FE_OFN1739_acc_fir_data_in_12_;
   wire FE_OFN1738_acc_fir_data_in_12_;
   wire FE_OFN1737_acc_fir_data_in_12_;
   wire FE_OFN1736_acc_fir_data_in_12_;
   wire FE_OFN1735_acc_fir_data_in_13_;
   wire FE_OFN1734_acc_fir_data_in_13_;
   wire FE_OFN1733_acc_fir_data_in_13_;
   wire FE_OFN1732_acc_fir_data_in_13_;
   wire FE_OFN1731_acc_fir_data_in_13_;
   wire FE_OFN1730_acc_fir_data_in_14_;
   wire FE_OFN1729_acc_fir_data_in_14_;
   wire FE_OFN1728_acc_fir_data_in_14_;
   wire FE_OFN1727_acc_fir_data_in_14_;
   wire FE_OFN1726_acc_fir_data_in_14_;
   wire FE_OFN1725_acc_fir_data_in_14_;
   wire FE_OFN1724_acc_fir_data_in_14_;
   wire FE_OFN1723_acc_fir_data_in_15_;
   wire FE_OFN1722_acc_fir_data_in_15_;
   wire FE_OFN1721_acc_fir_data_in_15_;
   wire FE_OFN1720_acc_fir_data_in_15_;
   wire FE_OFN1719_acc_fir_data_in_15_;
   wire FE_OFN1718_acc_fir_data_in_16_;
   wire FE_OFN1717_acc_fir_data_in_16_;
   wire FE_OFN1716_acc_fir_data_in_16_;
   wire FE_OFN1715_acc_fir_data_in_16_;
   wire FE_OFN1714_acc_fir_data_in_16_;
   wire FE_OFN1713_acc_fir_data_in_16_;
   wire FE_OFN1712_acc_fir_data_in_16_;
   wire FE_OFN1711_acc_fir_data_in_17_;
   wire FE_OFN1710_acc_fir_data_in_17_;
   wire FE_OFN1709_acc_fir_data_in_17_;
   wire FE_OFN1708_acc_fir_data_in_17_;
   wire FE_OFN1707_acc_fir_data_in_17_;
   wire FE_OFN1706_acc_fir_data_in_18_;
   wire FE_OFN1705_acc_fir_data_in_18_;
   wire FE_OFN1704_acc_fir_data_in_18_;
   wire FE_OFN1703_acc_fir_data_in_18_;
   wire FE_OFN1702_acc_fir_data_in_18_;
   wire FE_OFN1701_acc_fir_data_in_19_;
   wire FE_OFN1700_acc_fir_data_in_19_;
   wire FE_OFN1699_acc_fir_data_in_19_;
   wire FE_OFN1698_acc_fir_data_in_19_;
   wire FE_OFN1697_acc_fir_data_in_19_;
   wire FE_OFN1696_acc_fir_data_in_19_;
   wire FE_OFN1695_acc_fir_data_in_19_;
   wire FE_OFN1694_acc_fir_data_in_20_;
   wire FE_OFN1693_acc_fir_data_in_20_;
   wire FE_OFN1692_acc_fir_data_in_20_;
   wire FE_OFN1691_acc_fir_data_in_20_;
   wire FE_OFN1690_acc_fir_data_in_20_;
   wire FE_OFN1689_acc_fir_data_in_21_;
   wire FE_OFN1688_acc_fir_data_in_21_;
   wire FE_OFN1687_acc_fir_data_in_21_;
   wire FE_OFN1686_acc_fir_data_in_21_;
   wire FE_OFN1685_acc_fir_data_in_21_;
   wire FE_OFN1684_acc_fir_data_in_21_;
   wire FE_OFN1683_acc_fir_data_in_21_;
   wire FE_OFN1682_acc_fir_data_in_22_;
   wire FE_OFN1681_acc_fir_data_in_22_;
   wire FE_OFN1680_acc_fir_data_in_22_;
   wire FE_OFN1679_acc_fir_data_in_22_;
   wire FE_OFN1678_acc_fir_data_in_22_;
   wire FE_OFN1677_acc_fir_data_in_23_;
   wire FE_OFN1676_acc_fir_data_in_23_;
   wire FE_OFN1675_acc_fir_data_in_23_;
   wire FE_OFN1674_acc_fir_data_in_23_;
   wire FE_OFN1673_acc_fir_data_in_23_;
   wire FE_OFN1672_acc_fir_data_in_23_;
   wire FE_OFN1671_acc_fir_data_in_23_;
   wire FE_OFN1670_acc_fir_data_in_24_;
   wire FE_OFN1669_acc_fir_data_in_24_;
   wire FE_OFN1668_acc_fir_data_in_24_;
   wire FE_OFN1667_acc_fir_data_in_24_;
   wire FE_OFN1666_acc_fir_data_in_24_;
   wire FE_OFN1665_acc_fir_data_in_25_;
   wire FE_OFN1664_acc_fir_data_in_25_;
   wire FE_OFN1663_acc_fir_data_in_25_;
   wire FE_OFN1662_acc_fir_data_in_25_;
   wire FE_OFN1661_acc_fir_data_in_25_;
   wire FE_OFN1660_acc_fir_data_in_26_;
   wire FE_OFN1659_acc_fir_data_in_26_;
   wire FE_OFN1658_acc_fir_data_in_26_;
   wire FE_OFN1657_acc_fir_data_in_26_;
   wire FE_OFN1656_acc_fir_data_in_26_;
   wire FE_OFN1655_acc_fir_data_in_27_;
   wire FE_OFN1654_acc_fir_data_in_27_;
   wire FE_OFN1653_acc_fir_data_in_27_;
   wire FE_OFN1652_acc_fir_data_in_27_;
   wire FE_OFN1651_acc_fir_data_in_27_;
   wire FE_OFN1650_acc_fir_data_in_28_;
   wire FE_OFN1649_acc_fir_data_in_28_;
   wire FE_OFN1648_acc_fir_data_in_28_;
   wire FE_OFN1647_acc_fir_data_in_28_;
   wire FE_OFN1646_acc_fir_data_in_28_;
   wire FE_OFN1645_acc_fir_data_in_29_;
   wire FE_OFN1644_acc_fir_data_in_29_;
   wire FE_OFN1643_acc_fir_data_in_29_;
   wire FE_OFN1642_acc_fir_data_in_29_;
   wire FE_OFN1641_acc_fir_data_in_29_;
   wire FE_OFN1640_acc_fir_data_in_29_;
   wire FE_OFN1639_acc_fir_data_in_29_;
   wire FE_OFN1638_acc_fir_data_in_29_;
   wire FE_OFN1637_acc_fir_data_in_30_;
   wire FE_OFN1636_acc_fir_data_in_30_;
   wire FE_OFN1635_acc_fir_data_in_30_;
   wire FE_OFN1634_acc_fir_data_in_30_;
   wire FE_OFN1633_acc_fir_data_in_30_;
   wire FE_OFN1632_acc_fir_data_in_31_;
   wire FE_OFN1631_acc_fir_data_in_31_;
   wire FE_OFN1630_acc_fir_data_in_31_;
   wire FE_OFN1629_acc_fir_data_in_31_;
   wire FE_OFN1628_acc_fir_data_in_31_;
   wire FE_OFN1627_acc_fft_data_in_0_;
   wire FE_OFN1626_acc_fft_data_in_0_;
   wire FE_OFN1625_acc_fft_data_in_0_;
   wire FE_OFN1624_acc_fft_data_in_0_;
   wire FE_OFN1623_acc_fft_data_in_0_;
   wire FE_OFN1622_acc_fft_data_in_0_;
   wire FE_OFN1621_acc_fft_data_in_1_;
   wire FE_OFN1620_acc_fft_data_in_1_;
   wire FE_OFN1619_acc_fft_data_in_1_;
   wire FE_OFN1618_acc_fft_data_in_1_;
   wire FE_OFN1617_acc_fft_data_in_1_;
   wire FE_OFN1616_acc_fft_data_in_1_;
   wire FE_OFN1615_acc_fft_data_in_1_;
   wire FE_OFN1614_acc_fft_data_in_2_;
   wire FE_OFN1613_acc_fft_data_in_2_;
   wire FE_OFN1612_acc_fft_data_in_2_;
   wire FE_OFN1611_acc_fft_data_in_2_;
   wire FE_OFN1610_acc_fft_data_in_2_;
   wire FE_OFN1609_acc_fft_data_in_2_;
   wire FE_OFN1608_acc_fft_data_in_2_;
   wire FE_OFN1607_acc_fft_data_in_3_;
   wire FE_OFN1606_acc_fft_data_in_3_;
   wire FE_OFN1605_acc_fft_data_in_3_;
   wire FE_OFN1604_acc_fft_data_in_3_;
   wire FE_OFN1603_acc_fft_data_in_3_;
   wire FE_OFN1602_acc_fft_data_in_4_;
   wire FE_OFN1601_acc_fft_data_in_4_;
   wire FE_OFN1600_acc_fft_data_in_4_;
   wire FE_OFN1599_acc_fft_data_in_4_;
   wire FE_OFN1598_acc_fft_data_in_4_;
   wire FE_OFN1597_acc_fft_data_in_4_;
   wire FE_OFN1596_acc_fft_data_in_4_;
   wire FE_OFN1595_acc_fft_data_in_5_;
   wire FE_OFN1594_acc_fft_data_in_5_;
   wire FE_OFN1593_acc_fft_data_in_5_;
   wire FE_OFN1592_acc_fft_data_in_5_;
   wire FE_OFN1591_acc_fft_data_in_5_;
   wire FE_OFN1590_acc_fft_data_in_6_;
   wire FE_OFN1589_acc_fft_data_in_6_;
   wire FE_OFN1588_acc_fft_data_in_6_;
   wire FE_OFN1587_acc_fft_data_in_6_;
   wire FE_OFN1586_acc_fft_data_in_6_;
   wire FE_OFN1585_acc_fft_data_in_6_;
   wire FE_OFN1584_acc_fft_data_in_7_;
   wire FE_OFN1583_acc_fft_data_in_7_;
   wire FE_OFN1582_acc_fft_data_in_7_;
   wire FE_OFN1581_acc_fft_data_in_7_;
   wire FE_OFN1580_acc_fft_data_in_7_;
   wire FE_OFN1579_acc_fft_data_in_8_;
   wire FE_OFN1578_acc_fft_data_in_8_;
   wire FE_OFN1577_acc_fft_data_in_8_;
   wire FE_OFN1576_acc_fft_data_in_8_;
   wire FE_OFN1575_acc_fft_data_in_8_;
   wire FE_OFN1574_acc_fft_data_in_8_;
   wire FE_OFN1573_acc_fft_data_in_9_;
   wire FE_OFN1572_acc_fft_data_in_9_;
   wire FE_OFN1571_acc_fft_data_in_9_;
   wire FE_OFN1570_acc_fft_data_in_9_;
   wire FE_OFN1569_acc_fft_data_in_9_;
   wire FE_OFN1568_acc_fft_data_in_10_;
   wire FE_OFN1567_acc_fft_data_in_10_;
   wire FE_OFN1566_acc_fft_data_in_10_;
   wire FE_OFN1565_acc_fft_data_in_10_;
   wire FE_OFN1564_acc_fft_data_in_10_;
   wire FE_OFN1563_acc_fft_data_in_11_;
   wire FE_OFN1562_acc_fft_data_in_11_;
   wire FE_OFN1561_acc_fft_data_in_11_;
   wire FE_OFN1560_acc_fft_data_in_11_;
   wire FE_OFN1559_acc_fft_data_in_11_;
   wire FE_OFN1558_acc_fft_data_in_12_;
   wire FE_OFN1557_acc_fft_data_in_12_;
   wire FE_OFN1556_acc_fft_data_in_12_;
   wire FE_OFN1555_acc_fft_data_in_12_;
   wire FE_OFN1554_acc_fft_data_in_12_;
   wire FE_OFN1553_acc_fft_data_in_12_;
   wire FE_OFN1552_acc_fft_data_in_13_;
   wire FE_OFN1551_acc_fft_data_in_13_;
   wire FE_OFN1550_acc_fft_data_in_13_;
   wire FE_OFN1549_acc_fft_data_in_13_;
   wire FE_OFN1548_acc_fft_data_in_13_;
   wire FE_OFN1547_acc_fft_data_in_14_;
   wire FE_OFN1546_acc_fft_data_in_14_;
   wire FE_OFN1545_acc_fft_data_in_14_;
   wire FE_OFN1544_acc_fft_data_in_14_;
   wire FE_OFN1543_acc_fft_data_in_14_;
   wire FE_OFN1542_acc_fft_data_in_15_;
   wire FE_OFN1541_acc_fft_data_in_15_;
   wire FE_OFN1540_acc_fft_data_in_15_;
   wire FE_OFN1539_acc_fft_data_in_15_;
   wire FE_OFN1538_acc_fft_data_in_15_;
   wire FE_OFN1537_acc_fft_data_in_16_;
   wire FE_OFN1536_acc_fft_data_in_16_;
   wire FE_OFN1535_acc_fft_data_in_16_;
   wire FE_OFN1534_acc_fft_data_in_16_;
   wire FE_OFN1533_acc_fft_data_in_16_;
   wire FE_OFN1532_acc_fft_data_in_17_;
   wire FE_OFN1531_acc_fft_data_in_17_;
   wire FE_OFN1530_acc_fft_data_in_17_;
   wire FE_OFN1529_acc_fft_data_in_17_;
   wire FE_OFN1528_acc_fft_data_in_17_;
   wire FE_OFN1527_acc_fft_data_in_17_;
   wire FE_OFN1526_acc_fft_data_in_18_;
   wire FE_OFN1525_acc_fft_data_in_18_;
   wire FE_OFN1524_acc_fft_data_in_18_;
   wire FE_OFN1523_acc_fft_data_in_18_;
   wire FE_OFN1522_acc_fft_data_in_18_;
   wire FE_OFN1521_acc_fft_data_in_18_;
   wire FE_OFN1520_acc_fft_data_in_18_;
   wire FE_OFN1519_acc_fft_data_in_19_;
   wire FE_OFN1518_acc_fft_data_in_19_;
   wire FE_OFN1517_acc_fft_data_in_19_;
   wire FE_OFN1516_acc_fft_data_in_19_;
   wire FE_OFN1515_acc_fft_data_in_19_;
   wire FE_OFN1514_acc_fft_data_in_20_;
   wire FE_OFN1513_acc_fft_data_in_20_;
   wire FE_OFN1512_acc_fft_data_in_20_;
   wire FE_OFN1511_acc_fft_data_in_20_;
   wire FE_OFN1510_acc_fft_data_in_20_;
   wire FE_OFN1509_acc_fft_data_in_21_;
   wire FE_OFN1508_acc_fft_data_in_21_;
   wire FE_OFN1507_acc_fft_data_in_21_;
   wire FE_OFN1506_acc_fft_data_in_21_;
   wire FE_OFN1505_acc_fft_data_in_21_;
   wire FE_OFN1504_acc_fft_data_in_22_;
   wire FE_OFN1503_acc_fft_data_in_22_;
   wire FE_OFN1502_acc_fft_data_in_22_;
   wire FE_OFN1501_acc_fft_data_in_22_;
   wire FE_OFN1500_acc_fft_data_in_22_;
   wire FE_OFN1499_acc_fft_data_in_22_;
   wire FE_OFN1498_acc_fft_data_in_22_;
   wire FE_OFN1497_acc_fft_data_in_23_;
   wire FE_OFN1496_acc_fft_data_in_23_;
   wire FE_OFN1495_acc_fft_data_in_23_;
   wire FE_OFN1494_acc_fft_data_in_23_;
   wire FE_OFN1493_acc_fft_data_in_23_;
   wire FE_OFN1492_acc_fft_data_in_24_;
   wire FE_OFN1491_acc_fft_data_in_24_;
   wire FE_OFN1490_acc_fft_data_in_24_;
   wire FE_OFN1489_acc_fft_data_in_24_;
   wire FE_OFN1488_acc_fft_data_in_24_;
   wire FE_OFN1487_acc_fft_data_in_25_;
   wire FE_OFN1486_acc_fft_data_in_25_;
   wire FE_OFN1485_acc_fft_data_in_25_;
   wire FE_OFN1484_acc_fft_data_in_25_;
   wire FE_OFN1483_acc_fft_data_in_25_;
   wire FE_OFN1482_acc_fft_data_in_26_;
   wire FE_OFN1481_acc_fft_data_in_26_;
   wire FE_OFN1480_acc_fft_data_in_26_;
   wire FE_OFN1479_acc_fft_data_in_26_;
   wire FE_OFN1478_acc_fft_data_in_26_;
   wire FE_OFN1477_acc_fft_data_in_27_;
   wire FE_OFN1476_acc_fft_data_in_27_;
   wire FE_OFN1475_acc_fft_data_in_27_;
   wire FE_OFN1474_acc_fft_data_in_27_;
   wire FE_OFN1473_acc_fft_data_in_27_;
   wire FE_OFN1472_acc_fft_data_in_28_;
   wire FE_OFN1471_acc_fft_data_in_28_;
   wire FE_OFN1470_acc_fft_data_in_28_;
   wire FE_OFN1469_acc_fft_data_in_28_;
   wire FE_OFN1468_acc_fft_data_in_28_;
   wire FE_OFN1467_acc_fft_data_in_29_;
   wire FE_OFN1466_acc_fft_data_in_29_;
   wire FE_OFN1465_acc_fft_data_in_29_;
   wire FE_OFN1464_acc_fft_data_in_29_;
   wire FE_OFN1463_acc_fft_data_in_29_;
   wire FE_OFN1462_acc_fft_data_in_30_;
   wire FE_OFN1461_acc_fft_data_in_30_;
   wire FE_OFN1460_acc_fft_data_in_30_;
   wire FE_OFN1459_acc_fft_data_in_30_;
   wire FE_OFN1458_acc_fft_data_in_30_;
   wire FE_OFN1457_acc_fft_data_in_31_;
   wire FE_OFN1456_acc_fft_data_in_31_;
   wire FE_OFN1455_acc_fft_data_in_31_;
   wire FE_OFN1454_acc_fft_data_in_31_;
   wire FE_OFN1453_acc_fft_data_in_31_;
   wire FE_OFN1452_acc_fft_data_in_31_;
   wire FE_OFN1451_acc_fir_put;
   wire FE_OFN1450_acc_fir_get;
   wire FE_OFN1449_acc_fft_put;
   wire FE_OFN1448_acc_fft_get;
   wire FE_OFN1447_reset;
   wire FE_OFN1446_router_addr_calc_fir_read_calc_count_0_;
   wire FE_OFN1445_router_addr_calc_fir_write_calc_count_0_;
   wire FE_OFN1444_router_addr_calc_fft_read_calc_count_0_;
   wire FE_OFN1443_router_addr_calc_fft_write_calc_count_0_;
   wire FE_OFN1442_router_addr_calc_iir_write_calc_count_0_;
   wire FE_OFN1441_router_addr_calc_iir_write_calc_count_16_;
   wire FE_OFN1440_router_addr_calc_iir_write_calc_count_19_;
   wire FE_OFN1439_router_addr_calc_iir_write_calc_count_27_;
   wire FE_OFN1438_router_data_from_fft;
   wire FE_OFN1437_n8093;
   wire FE_OFN1436_n8093;
   wire FE_OFN1435_n8093;
   wire FE_OFN1434_n8093;
   wire FE_OFN1433_n8093;
   wire FE_OFN1432_n8092;
   wire FE_OFN1431_n8092;
   wire FE_OFN1430_n8092;
   wire FE_OFN1429_n8092;
   wire FE_OFN1428_n8091;
   wire FE_OFN1427_n8091;
   wire FE_OFN1426_n8091;
   wire FE_OFN1425_n8091;
   wire FE_OFN1424_n8090;
   wire FE_OFN1423_n8090;
   wire FE_OFN1422_n8090;
   wire FE_OFN1421_n8090;
   wire FE_OFN1420_n8090;
   wire FE_OFN1419_n8089;
   wire FE_OFN1418_n8089;
   wire FE_OFN1417_n8089;
   wire FE_OFN1416_n8089;
   wire FE_OFN1415_n8088;
   wire FE_OFN1414_n8088;
   wire FE_OFN1413_n8088;
   wire FE_OFN1412_n8088;
   wire FE_OFN1411_n8087;
   wire FE_OFN1410_n8087;
   wire FE_OFN1409_n8087;
   wire FE_OFN1408_n8087;
   wire FE_OFN1407_n8087;
   wire FE_OFN1406_n8086;
   wire FE_OFN1405_n8086;
   wire FE_OFN1404_n8086;
   wire FE_OFN1403_n8086;
   wire FE_OFN1402_n8085;
   wire FE_OFN1401_n8085;
   wire FE_OFN1400_n8085;
   wire FE_OFN1399_n8085;
   wire FE_OFN1398_n8084;
   wire FE_OFN1397_n8084;
   wire FE_OFN1396_n8084;
   wire FE_OFN1395_n8084;
   wire FE_OFN1394_n8084;
   wire FE_OFN1393_n8083;
   wire FE_OFN1392_n8083;
   wire FE_OFN1391_n8083;
   wire FE_OFN1390_n8083;
   wire FE_OFN1389_n8083;
   wire FE_OFN1388_n8082;
   wire FE_OFN1387_n8082;
   wire FE_OFN1386_n8082;
   wire FE_OFN1385_n8082;
   wire FE_OFN1384_n8082;
   wire FE_OFN1383_n8081;
   wire FE_OFN1382_n8081;
   wire FE_OFN1381_n8081;
   wire FE_OFN1380_n8081;
   wire FE_OFN1379_n8080;
   wire FE_OFN1378_n8080;
   wire FE_OFN1377_n8080;
   wire FE_OFN1376_n8080;
   wire FE_OFN1375_n8078;
   wire FE_OFN1374_n8078;
   wire FE_OFN1373_n8078;
   wire FE_OFN1372_n8078;
   wire FE_OFN1371_n8078;
   wire FE_OFN1370_n8077;
   wire FE_OFN1369_n8077;
   wire FE_OFN1368_n8077;
   wire FE_OFN1367_n8077;
   wire FE_OFN1366_n8077;
   wire FE_OFN1365_n8076;
   wire FE_OFN1364_n8076;
   wire FE_OFN1363_n8076;
   wire FE_OFN1362_n8076;
   wire FE_OFN1361_n8075;
   wire FE_OFN1360_n8075;
   wire FE_OFN1359_n8075;
   wire FE_OFN1358_n8075;
   wire FE_OFN1357_n8075;
   wire FE_OFN1356_n8074;
   wire FE_OFN1355_n8074;
   wire FE_OFN1354_n8074;
   wire FE_OFN1353_n8074;
   wire FE_OFN1352_n8073;
   wire FE_OFN1351_n8073;
   wire FE_OFN1350_n8073;
   wire FE_OFN1349_n8073;
   wire FE_OFN1348_n8072;
   wire FE_OFN1347_n8072;
   wire FE_OFN1346_n8072;
   wire FE_OFN1345_n8072;
   wire FE_OFN1344_n8072;
   wire FE_OFN1343_n8071;
   wire FE_OFN1342_n8071;
   wire FE_OFN1341_n8071;
   wire FE_OFN1340_n8071;
   wire FE_OFN1339_n8071;
   wire FE_OFN1338_n8070;
   wire FE_OFN1337_n8070;
   wire FE_OFN1336_n8070;
   wire FE_OFN1335_n8070;
   wire FE_OFN1334_n8069;
   wire FE_OFN1333_n8069;
   wire FE_OFN1332_n8069;
   wire FE_OFN1331_n8069;
   wire FE_OFN1330_n8068;
   wire FE_OFN1329_n8068;
   wire FE_OFN1328_n8068;
   wire FE_OFN1327_n8068;
   wire FE_OFN1326_n8067;
   wire FE_OFN1325_n8067;
   wire FE_OFN1324_n8067;
   wire FE_OFN1323_n8067;
   wire FE_OFN1322_n8066;
   wire FE_OFN1321_n8066;
   wire FE_OFN1320_n8066;
   wire FE_OFN1319_n8066;
   wire FE_OFN1318_n8066;
   wire FE_OFN1317_n8065;
   wire FE_OFN1316_n8065;
   wire FE_OFN1315_n8065;
   wire FE_OFN1314_n8065;
   wire FE_OFN1313_n8094;
   wire FE_OFN1312_n8094;
   wire FE_OFN1311_n8094;
   wire FE_OFN1310_n8094;
   wire FE_OFN1309_n8079;
   wire FE_OFN1308_n8079;
   wire FE_OFN1307_n8079;
   wire FE_OFN1306_n8079;
   wire FE_OFN1305_n8060;
   wire FE_OFN1304_n8060;
   wire FE_OFN1303_n8060;
   wire FE_OFN1302_n8060;
   wire FE_OFN1301_n8060;
   wire FE_OFN1300_iir_enable;
   wire FE_OFN1299_iir_enable;
   wire FE_OFN1298_iir_enable;
   wire FE_OFN1297_iir_enable;
   wire FE_OFN1296_iir_enable;
   wire FE_OFN1295_iir_enable;
   wire FE_OFN1294_iir_enable;
   wire FE_OFN1293_iir_enable;
   wire FE_OFN1292_iir_enable;
   wire FE_OFN1291_iir_enable;
   wire FE_OFN1290_iir_enable;
   wire FE_OFN1289_iir_enable;
   wire FE_OFN1288_iir_enable;
   wire FE_OFN1287_iir_enable;
   wire FE_OFN1286_iir_enable;
   wire FE_OFN1285_router_ram_read_enable_reg;
   wire FE_OFN1284_router_ram_read_enable_reg;
   wire FE_OFN1283_router_fft_write_done;
   wire FE_OFN1282_router_fft_get_req_reg;
   wire FE_OFN1281_router_addr_calc_iir_write_calc_count_5_;
   wire FE_OFN1280_router_addr_calc_iir_write_calc_count_9_;
   wire FE_OFN1279_n7328;
   wire FE_OFN1278_n7333;
   wire FE_OFN1277_n7308;
   wire FE_OFN1276_router_addr_calc_fir_read_calc_count_5_;
   wire FE_OFN1275_n7353;
   wire FE_OFN1274_n7358;
   wire FE_OFN1273_router_addr_calc_fft_read_calc_count_5_;
   wire FE_OFN1272_router_addr_calc_fir_write_calc_count_5_;
   wire FE_OFN1271_router_addr_calc_fir_read_calc_count_15_;
   wire FE_OFN1270_router_addr_calc_fft_write_calc_count_15_;
   wire FE_OFN1269_router_addr_calc_fir_read_calc_count_9_;
   wire FE_OFN1268_router_addr_calc_fft_write_calc_count_9_;
   wire FE_OFN1267_router_addr_calc_fft_read_calc_count_9_;
   wire FE_OFN1266_router_addr_calc_fir_write_calc_count_9_;
   wire FE_OFN1265_n7303;
   wire FE_OFN1264_router_addr_calc_fir_write_calc_count_16_;
   wire FE_OFN1263_router_addr_calc_fft_read_calc_count_16_;
   wire FE_OFN1262_n7298;
   wire FE_OFN1261_router_addr_calc_fir_write_calc_count_19_;
   wire FE_OFN1260_router_addr_calc_fir_read_calc_count_19_;
   wire FE_OFN1259_router_addr_calc_fft_write_calc_count_19_;
   wire FE_OFN1258_router_addr_calc_fft_read_calc_count_19_;
   wire FE_OFN1257_n7165;
   wire FE_OFN1256_n7288;
   wire FE_OFN1255_n7402;
   wire FE_OFN1254_n7159;
   wire FE_OFN1253_n7283;
   wire FE_OFN1252_n7397;
   wire FE_OFN1251_n7153;
   wire FE_OFN1250_n7278;
   wire FE_OFN1249_n7392;
   wire FE_OFN1248_router_addr_calc_fir_write_calc_count_23_;
   wire FE_OFN1247_router_addr_calc_fir_read_calc_count_23_;
   wire FE_OFN1246_router_addr_calc_fft_write_calc_count_23_;
   wire FE_OFN1245_router_addr_calc_fft_read_calc_count_23_;
   wire FE_OFN1244_router_addr_calc_iir_write_calc_count_23_;
   wire FE_OFN1243_n7273;
   wire FE_OFN1242_n7268;
   wire FE_OFN1241_n7264;
   wire FE_OFN1240_router_addr_calc_fir_write_calc_count_27_;
   wire FE_OFN1239_router_addr_calc_fir_read_calc_count_27_;
   wire FE_OFN1238_router_addr_calc_fft_write_calc_count_27_;
   wire FE_OFN1237_router_addr_calc_fft_read_calc_count_27_;
   wire FE_OFN1236_n7259;
   wire FE_OFN1235_n7254;
   wire FE_OFN1234_n7492;
   wire FE_OFN1233_router_addr_calc_fft_write_calc_count_29_;
   wire FE_OFN1232_n7368;
   wire FE_OFN1231_router_addr_calc_fir_write_calc_count_30_;
   wire FE_OFN1230_router_addr_calc_fir_read_calc_count_30_;
   wire FE_OFN1229_router_addr_calc_fft_read_calc_count_30_;
   wire FE_OFN1228_router_addr_calc_fft_write_calc_count_31_;
   wire FE_OFN1227_n8063;
   wire FE_OFN1226_n8063;
   wire FE_OFN1225_n8063;
   wire FE_OFN1224_n8063;
   wire FE_OFN1223_n8063;
   wire FE_OFN1222_n8064;
   wire FE_OFN1221_n8064;
   wire FE_OFN1220_n8064;
   wire FE_OFN1219_n8064;
   wire FE_OFN1218_n8064;
   wire FE_OFN1217_n3478;
   wire FE_OFN1216_n8061;
   wire FE_OFN1215_n8061;
   wire FE_OFN1214_n8061;
   wire FE_OFN1213_n8061;
   wire FE_OFN1212_n8061;
   wire FE_OFN1211_n8062;
   wire FE_OFN1210_n8062;
   wire FE_OFN1209_n8062;
   wire FE_OFN1208_n8062;
   wire FE_OFN1207_router_addr_calc_iir_write_calc_counter_N212;
   wire FE_OFN1206_router_addr_calc_iir_write_calc_counter_N212;
   wire FE_OFN1205_router_addr_calc_iir_write_calc_counter_N212;
   wire FE_OFN1204_router_addr_calc_iir_write_calc_counter_N212;
   wire FE_OFN1203_router_addr_calc_iir_write_calc_counter_N212;
   wire FE_OFN1202_router_addr_calc_iir_write_calc_counter_N212;
   wire FE_OFN1201_router_addr_calc_iir_write_calc_counter_N212;
   wire FE_OFN1200_router_addr_calc_iir_write_calc_counter_N212;
   wire FE_OFN1199_router_addr_calc_iir_write_calc_counter_N212;
   wire FE_OFN1198_n7023;
   wire FE_OFN1197_n7023;
   wire FE_OFN1196_n7023;
   wire FE_OFN1195_n7023;
   wire FE_OFN1194_n7023;
   wire FE_OFN1193_n7023;
   wire FE_OFN1192_n7022;
   wire FE_OFN1191_n7022;
   wire FE_OFN1190_n7022;
   wire FE_OFN1189_n7020;
   wire FE_OFN1188_n7020;
   wire FE_OFN1187_n7020;
   wire FE_OFN1186_n7020;
   wire FE_OFN1185_n7020;
   wire FE_OFN1184_n7020;
   wire FE_OFN1183_n7020;
   wire FE_OFN1182_n7020;
   wire FE_OFN1181_n7020;
   wire FE_OFN1180_n7020;
   wire FE_OFN1179_n7020;
   wire FE_OFN1178_n7021;
   wire FE_OFN1177_n7021;
   wire FE_OFN1176_n7021;
   wire FE_OFN1175_n7021;
   wire FE_OFN1174_n7021;
   wire FE_OFN1173_n7021;
   wire FE_OFN1172_n7021;
   wire FE_OFN1171_n7021;
   wire FE_OFN1170_n7021;
   wire FE_OFN1169_n7021;
   wire FE_OFN1168_n7021;
   wire FE_OFN1167_n7019;
   wire FE_OFN1166_n7019;
   wire FE_OFN1165_n7019;
   wire FE_OFN1164_n7019;
   wire FE_OFN1163_n7019;
   wire FE_OFN1162_n7019;
   wire FE_OFN1161_n7019;
   wire FE_OFN1160_n7019;
   wire FE_OFN1159_n7019;
   wire FE_OFN1158_n7019;
   wire FE_OFN1157_n1609;
   wire FE_OFN1156_n1609;
   wire FE_OFN1155_n1609;
   wire FE_OFN1154_n1609;
   wire FE_OFN1153_n1609;
   wire FE_OFN1152_n1609;
   wire FE_OFN1151_n1609;
   wire FE_OFN1150_n1609;
   wire FE_OFN1149_n1609;
   wire FE_OFN1148_n1609;
   wire FE_OFN1147_n585;
   wire FE_OFN1146_n585;
   wire FE_OFN1145_n585;
   wire FE_OFN1144_n585;
   wire FE_OFN1143_n585;
   wire FE_OFN1142_n585;
   wire FE_OFN1141_n585;
   wire FE_OFN1140_n585;
   wire FE_OFN1139_n585;
   wire FE_OFN1138_n585;
   wire FE_OFN1137_n2505;
   wire FE_OFN1136_n2505;
   wire FE_OFN1135_n2505;
   wire FE_OFN1134_n2505;
   wire FE_OFN1133_n2505;
   wire FE_OFN1132_n2441;
   wire FE_OFN1131_n2441;
   wire FE_OFN1130_n2441;
   wire FE_OFN1129_n2441;
   wire FE_OFN1128_n2377;
   wire FE_OFN1127_n2377;
   wire FE_OFN1126_n2377;
   wire FE_OFN1125_n2377;
   wire FE_OFN1124_n2377;
   wire FE_OFN1123_n2313;
   wire FE_OFN1122_n2313;
   wire FE_OFN1121_n2313;
   wire FE_OFN1120_n2313;
   wire FE_OFN1119_n2249;
   wire FE_OFN1118_n2249;
   wire FE_OFN1117_n2249;
   wire FE_OFN1116_n2249;
   wire FE_OFN1115_n2249;
   wire FE_OFN1114_n2185;
   wire FE_OFN1113_n2185;
   wire FE_OFN1112_n2185;
   wire FE_OFN1111_n2185;
   wire FE_OFN1110_n2121;
   wire FE_OFN1109_n2121;
   wire FE_OFN1108_n2121;
   wire FE_OFN1107_n2121;
   wire FE_OFN1106_n2121;
   wire FE_OFN1105_n2057;
   wire FE_OFN1104_n2057;
   wire FE_OFN1103_n2057;
   wire FE_OFN1102_n2057;
   wire FE_OFN1101_n1993;
   wire FE_OFN1100_n1993;
   wire FE_OFN1099_n1993;
   wire FE_OFN1098_n1993;
   wire FE_OFN1097_n1993;
   wire FE_OFN1096_n1929;
   wire FE_OFN1095_n1929;
   wire FE_OFN1094_n1929;
   wire FE_OFN1093_n1929;
   wire FE_OFN1092_n1865;
   wire FE_OFN1091_n1865;
   wire FE_OFN1090_n1865;
   wire FE_OFN1089_n1865;
   wire FE_OFN1088_n1801;
   wire FE_OFN1087_n1801;
   wire FE_OFN1086_n1801;
   wire FE_OFN1085_n1801;
   wire FE_OFN1084_n1737;
   wire FE_OFN1083_n1737;
   wire FE_OFN1082_n1737;
   wire FE_OFN1081_n1737;
   wire FE_OFN1080_n1673;
   wire FE_OFN1079_n1673;
   wire FE_OFN1078_n1673;
   wire FE_OFN1077_n1673;
   wire FE_OFN1076_n1481;
   wire FE_OFN1075_n1481;
   wire FE_OFN1074_n1481;
   wire FE_OFN1073_n1481;
   wire FE_OFN1072_n1417;
   wire FE_OFN1071_n1417;
   wire FE_OFN1070_n1417;
   wire FE_OFN1069_n1417;
   wire FE_OFN1068_n1353;
   wire FE_OFN1067_n1353;
   wire FE_OFN1066_n1353;
   wire FE_OFN1065_n1353;
   wire FE_OFN1064_n1289;
   wire FE_OFN1063_n1289;
   wire FE_OFN1062_n1289;
   wire FE_OFN1061_n1289;
   wire FE_OFN1060_n1225;
   wire FE_OFN1059_n1225;
   wire FE_OFN1058_n1225;
   wire FE_OFN1057_n1225;
   wire FE_OFN1056_n1225;
   wire FE_OFN1055_n1161;
   wire FE_OFN1054_n1161;
   wire FE_OFN1053_n1161;
   wire FE_OFN1052_n1161;
   wire FE_OFN1051_n1097;
   wire FE_OFN1050_n1097;
   wire FE_OFN1049_n1097;
   wire FE_OFN1048_n1097;
   wire FE_OFN1047_n1033;
   wire FE_OFN1046_n1033;
   wire FE_OFN1045_n1033;
   wire FE_OFN1044_n1033;
   wire FE_OFN1043_n1033;
   wire FE_OFN1042_n969;
   wire FE_OFN1041_n969;
   wire FE_OFN1040_n969;
   wire FE_OFN1039_n969;
   wire FE_OFN1038_n905;
   wire FE_OFN1037_n905;
   wire FE_OFN1036_n905;
   wire FE_OFN1035_n905;
   wire FE_OFN1034_n905;
   wire FE_OFN1033_n841;
   wire FE_OFN1032_n841;
   wire FE_OFN1031_n841;
   wire FE_OFN1030_n841;
   wire FE_OFN1029_n777;
   wire FE_OFN1028_n777;
   wire FE_OFN1027_n777;
   wire FE_OFN1026_n777;
   wire FE_OFN1025_n713;
   wire FE_OFN1024_n713;
   wire FE_OFN1023_n713;
   wire FE_OFN1022_n713;
   wire FE_OFN1021_n649;
   wire FE_OFN1020_n649;
   wire FE_OFN1019_n649;
   wire FE_OFN1018_n649;
   wire FE_OFN1017_n2569;
   wire FE_OFN1016_n2569;
   wire FE_OFN1015_n2569;
   wire FE_OFN1014_n2569;
   wire FE_OFN1013_n1545;
   wire FE_OFN1012_n1545;
   wire FE_OFN1011_n1545;
   wire FE_OFN1010_n1545;
   wire FE_OFN1009_n1545;
   wire FE_OFN1008_n137;
   wire FE_OFN1007_n137;
   wire FE_OFN1006_n137;
   wire FE_OFN1005_n137;
   wire FE_OFN1004_n137;
   wire FE_OFN1003_n521;
   wire FE_OFN1002_n521;
   wire FE_OFN1001_n521;
   wire FE_OFN1000_n521;
   wire FE_OFN999_n521;
   wire FE_OFN998_n521;
   wire FE_OFN997_n521;
   wire FE_OFN996_n521;
   wire FE_OFN995_n521;
   wire FE_OFN994_n521;
   wire FE_OFN993_n9431;
   wire FE_OFN992_n9431;
   wire FE_OFN991_n9431;
   wire FE_OFN990_n9431;
   wire FE_OFN989_n9431;
   wire FE_OFN988_n9431;
   wire FE_OFN987_n9431;
   wire FE_OFN986_n9431;
   wire FE_OFN985_n9431;
   wire FE_OFN984_n9462;
   wire FE_OFN983_n9462;
   wire FE_OFN982_n9462;
   wire FE_OFN981_n9462;
   wire FE_OFN980_n9462;
   wire FE_OFN979_n9462;
   wire FE_OFN978_n9462;
   wire FE_OFN977_n9462;
   wire FE_OFN976_n9462;
   wire FE_OFN975_n9462;
   wire FE_OFN974_n9462;
   wire FE_OFN973_n7207;
   wire FE_OFN972_n3618;
   wire FE_OFN971_n3618;
   wire FE_OFN970_n3618;
   wire FE_OFN969_n3618;
   wire FE_OFN968_n3618;
   wire FE_OFN967_n3618;
   wire FE_OFN966_n3618;
   wire FE_OFN965_n3618;
   wire FE_OFN964_n3618;
   wire FE_OFN963_n3618;
   wire FE_OFN962_n3618;
   wire FE_OFN961_n5467;
   wire FE_OFN960_n3619;
   wire FE_OFN959_n3619;
   wire FE_OFN958_n3619;
   wire FE_OFN957_n3619;
   wire FE_OFN956_n3619;
   wire FE_OFN955_n3619;
   wire FE_OFN954_n3619;
   wire FE_OFN953_n3619;
   wire FE_OFN952_n3619;
   wire FE_OFN951_n3619;
   wire FE_OFN950_n3486;
   wire FE_OFN949_n3486;
   wire FE_OFN948_n3486;
   wire FE_OFN947_n3486;
   wire FE_OFN946_n3486;
   wire FE_OFN945_n3486;
   wire FE_OFN944_n3486;
   wire FE_OFN943_n3486;
   wire FE_OFN942_n3486;
   wire FE_OFN941_n3486;
   wire FE_OFN940_n3486;
   wire FE_OFN939_n3487;
   wire FE_OFN938_n3487;
   wire FE_OFN937_n3487;
   wire FE_OFN936_n3487;
   wire FE_OFN935_n3487;
   wire FE_OFN934_n3487;
   wire FE_OFN933_n3487;
   wire FE_OFN932_n3487;
   wire FE_OFN931_n3487;
   wire FE_OFN930_n3487;
   wire FE_OFN929_n3574;
   wire FE_OFN928_n3574;
   wire FE_OFN927_n3574;
   wire FE_OFN926_n3574;
   wire FE_OFN925_n3574;
   wire FE_OFN924_n3574;
   wire FE_OFN923_n3574;
   wire FE_OFN922_n3574;
   wire FE_OFN921_n3574;
   wire FE_OFN920_n3574;
   wire FE_OFN919_n3574;
   wire FE_OFN918_n3575;
   wire FE_OFN917_n3575;
   wire FE_OFN916_n3575;
   wire FE_OFN915_n3575;
   wire FE_OFN914_n3575;
   wire FE_OFN913_n3575;
   wire FE_OFN912_n3575;
   wire FE_OFN911_n3575;
   wire FE_OFN910_n3575;
   wire FE_OFN909_n3575;
   wire FE_OFN908_n3530;
   wire FE_OFN907_n3530;
   wire FE_OFN906_n3530;
   wire FE_OFN905_n3530;
   wire FE_OFN904_n3530;
   wire FE_OFN903_n3530;
   wire FE_OFN902_n3530;
   wire FE_OFN901_n3530;
   wire FE_OFN900_n3530;
   wire FE_OFN899_n3530;
   wire FE_OFN898_n3530;
   wire FE_OFN897_n3531;
   wire FE_OFN896_n3531;
   wire FE_OFN895_n3531;
   wire FE_OFN894_n3531;
   wire FE_OFN893_n3531;
   wire FE_OFN892_n3531;
   wire FE_OFN891_n3531;
   wire FE_OFN890_n3531;
   wire FE_OFN889_n3531;
   wire FE_OFN888_n3531;
   wire FE_OFN887_n3662;
   wire FE_OFN886_n3662;
   wire FE_OFN885_n3662;
   wire FE_OFN884_n3662;
   wire FE_OFN883_n3662;
   wire FE_OFN882_n3662;
   wire FE_OFN881_n3662;
   wire FE_OFN880_n3662;
   wire FE_OFN879_n3662;
   wire FE_OFN878_n3662;
   wire FE_OFN877_n3662;
   wire FE_OFN876_n3663;
   wire FE_OFN875_n3663;
   wire FE_OFN874_n3663;
   wire FE_OFN873_n3663;
   wire FE_OFN872_n3663;
   wire FE_OFN871_n3663;
   wire FE_OFN870_n3663;
   wire FE_OFN869_n3663;
   wire FE_OFN868_n3663;
   wire FE_OFN867_n3663;
   wire FE_OFN866_n7015;
   wire FE_OFN865_n7015;
   wire FE_OFN864_n7015;
   wire FE_OFN863_n7015;
   wire FE_OFN862_n7015;
   wire FE_OFN861_n7017;
   wire FE_OFN860_n7017;
   wire FE_OFN859_n7017;
   wire FE_OFN858_n7017;
   wire FE_OFN857_n7017;
   wire FE_OFN856_n7018;
   wire FE_OFN855_n7018;
   wire FE_OFN854_n7018;
   wire FE_OFN853_n7018;
   wire FE_OFN852_n7016;
   wire FE_OFN851_n7016;
   wire FE_OFN850_n7016;
   wire FE_OFN849_n7016;
   wire FE_OFN848_ram_write_enable;
   wire FE_OFN847_n7619;
   wire FE_OFN846_n7619;
   wire FE_OFN845_n7619;
   wire FE_OFN844_n7619;
   wire FE_OFN843_n7619;
   wire FE_OFN842_n7619;
   wire FE_OFN841_n7619;
   wire FE_OFN840_n7619;
   wire FE_OFN839_n7619;
   wire FE_OFN838_n7619;
   wire FE_OFN837_n7619;
   wire FE_OFN836_n7619;
   wire FE_OFN835_n7619;
   wire FE_OFN834_n7619;
   wire FE_OFN833_n7619;
   wire FE_OFN832_n7619;
   wire FE_OFN831_n7619;
   wire FE_OFN830_n7619;
   wire FE_OFN829_n7619;
   wire FE_OFN828_n7619;
   wire FE_OFN827_n7619;
   wire FE_OFN826_n7619;
   wire FE_OFN825_n7619;
   wire FE_OFN824_n7619;
   wire FE_OFN823_n7619;
   wire FE_OFN822_n7619;
   wire FE_OFN821_n7619;
   wire FE_OFN820_n7619;
   wire FE_OFN819_n7619;
   wire FE_OFN818_n7619;
   wire FE_OFN817_n7619;
   wire FE_OFN816_n7619;
   wire FE_OFN815_n7619;
   wire FE_OFN814_n7619;
   wire FE_OFN813_n7619;
   wire FE_OFN812_n7619;
   wire FE_OFN811_n7619;
   wire FE_OFN810_n7619;
   wire FE_OFN809_n7619;
   wire FE_OFN808_n7619;
   wire FE_OFN807_n7619;
   wire FE_OFN806_n7619;
   wire FE_OFN805_n7619;
   wire FE_OFN804_n7619;
   wire FE_OFN803_n7619;
   wire FE_OFN802_n7619;
   wire FE_OFN801_n7619;
   wire FE_OFN800_n7619;
   wire FE_OFN799_n7619;
   wire FE_OFN798_n7619;
   wire FE_OFN797_n7619;
   wire FE_OFN796_n7619;
   wire FE_OFN795_n7619;
   wire FE_OFN794_n7619;
   wire FE_OFN793_n7619;
   wire FE_OFN792_n7619;
   wire FE_OFN791_n7619;
   wire FE_OFN790_n7619;
   wire FE_OFN789_n7619;
   wire FE_OFN788_n7619;
   wire FE_OFN787_n7619;
   wire FE_OFN786_n7619;
   wire FE_OFN785_n7619;
   wire FE_OFN784_n7619;
   wire FE_OFN783_n7619;
   wire FE_OFN782_n7619;
   wire FE_OFN781_n7619;
   wire FE_OFN780_n7619;
   wire FE_OFN779_n7619;
   wire FE_OFN778_n7619;
   wire FE_OFN777_n7619;
   wire FE_OFN776_n3829;
   wire FE_OFN775_n3720;
   wire FE_OFN774_n3720;
   wire FE_OFN773_n3720;
   wire FE_OFN772_n3720;
   wire FE_OFN771_n3720;
   wire FE_OFN770_n3720;
   wire FE_OFN769_n3720;
   wire FE_OFN768_n3720;
   wire FE_OFN767_n3720;
   wire FE_OFN766_n3720;
   wire FE_OFN765_n3720;
   wire FE_OFN764_n3721;
   wire FE_OFN763_n3721;
   wire FE_OFN762_n3721;
   wire FE_OFN761_n3721;
   wire FE_OFN760_n3721;
   wire FE_OFN759_n3721;
   wire FE_OFN758_n3721;
   wire FE_OFN757_n3721;
   wire FE_OFN756_n3721;
   wire FE_OFN755_n3721;
   wire FE_OFN754_n3722;
   wire FE_OFN753_n3722;
   wire FE_OFN752_n3722;
   wire FE_OFN751_n3722;
   wire FE_OFN750_n3722;
   wire FE_OFN749_n3722;
   wire FE_OFN748_n3722;
   wire FE_OFN747_n3722;
   wire FE_OFN746_n3722;
   wire FE_OFN745_n3722;
   wire FE_OFN744_n4829;
   wire FE_OFN743_n4829;
   wire FE_OFN742_n4829;
   wire FE_OFN741_n4829;
   wire FE_OFN740_n4829;
   wire FE_OFN739_n4829;
   wire FE_OFN738_n4829;
   wire FE_OFN737_n4829;
   wire FE_OFN736_n4829;
   wire FE_OFN735_n4829;
   wire FE_OFN734_n8057;
   wire FE_OFN733_n8057;
   wire FE_OFN732_n8057;
   wire FE_OFN731_n8058;
   wire FE_OFN730_n8058;
   wire FE_OFN729_n8058;
   wire FE_OFN728_n4643;
   wire FE_OFN727_n4643;
   wire FE_OFN726_n4643;
   wire FE_OFN725_n4643;
   wire FE_OFN724_n4643;
   wire FE_OFN723_n4643;
   wire FE_OFN722_n4643;
   wire FE_OFN721_n4643;
   wire FE_OFN720_n4643;
   wire FE_OFN719_n4643;
   wire FE_OFN718_n8051;
   wire FE_OFN717_n8051;
   wire FE_OFN716_n4207;
   wire FE_OFN715_n4207;
   wire FE_OFN714_n4207;
   wire FE_OFN713_n4207;
   wire FE_OFN712_n4207;
   wire FE_OFN711_n4207;
   wire FE_OFN710_n4207;
   wire FE_OFN709_n4207;
   wire FE_OFN708_n3959;
   wire FE_OFN707_n3959;
   wire FE_OFN706_n3959;
   wire FE_OFN705_n3959;
   wire FE_OFN704_n3959;
   wire FE_OFN703_n3959;
   wire FE_OFN702_n3959;
   wire FE_OFN701_n3959;
   wire FE_OFN700_n3959;
   wire FE_OFN699_n3959;
   wire FE_OFN698_n8052;
   wire FE_OFN697_n8052;
   wire FE_OFN696_n8052;
   wire FE_OFN695_n4134;
   wire FE_OFN694_n4134;
   wire FE_OFN693_n4134;
   wire FE_OFN692_n4134;
   wire FE_OFN691_n4134;
   wire FE_OFN690_n4134;
   wire FE_OFN689_n4134;
   wire FE_OFN688_n4134;
   wire FE_OFN687_n4134;
   wire FE_OFN686_n4134;
   wire FE_OFN685_n4134;
   wire FE_OFN684_n4134;
   wire FE_OFN683_n4134;
   wire FE_OFN682_n8050;
   wire FE_OFN681_n8050;
   wire FE_OFN680_n8050;
   wire FE_OFN679_n8050;
   wire FE_OFN678_n7295;
   wire FE_OFN677_n4759;
   wire FE_OFN676_n4759;
   wire FE_OFN675_n4759;
   wire FE_OFN674_n4759;
   wire FE_OFN673_n4759;
   wire FE_OFN672_n4759;
   wire FE_OFN671_n4759;
   wire FE_OFN670_n4759;
   wire FE_OFN669_n4759;
   wire FE_OFN668_n4759;
   wire FE_OFN667_n4759;
   wire FE_OFN666_n4759;
   wire FE_OFN665_n8053;
   wire FE_OFN664_n8053;
   wire FE_OFN663_n4747;
   wire FE_OFN662_n4747;
   wire FE_OFN661_n4747;
   wire FE_OFN660_n4747;
   wire FE_OFN659_n4747;
   wire FE_OFN658_n4747;
   wire FE_OFN657_n4747;
   wire FE_OFN656_n4747;
   wire FE_OFN655_n4747;
   wire FE_OFN654_n4747;
   wire FE_OFN653_n4747;
   wire FE_OFN652_n4747;
   wire FE_OFN651_n4741;
   wire FE_OFN650_n4741;
   wire FE_OFN649_n4741;
   wire FE_OFN648_n4741;
   wire FE_OFN647_n4741;
   wire FE_OFN646_n4741;
   wire FE_OFN645_n4741;
   wire FE_OFN644_n4741;
   wire FE_OFN643_n4741;
   wire FE_OFN642_n4741;
   wire FE_OFN641_n4741;
   wire FE_OFN640_n4741;
   wire FE_OFN639_n4742;
   wire FE_OFN638_n4742;
   wire FE_OFN637_n4742;
   wire FE_OFN636_n4742;
   wire FE_OFN635_n4742;
   wire FE_OFN634_n4742;
   wire FE_OFN633_n4742;
   wire FE_OFN632_n4742;
   wire FE_OFN631_n4742;
   wire FE_OFN630_n4742;
   wire FE_OFN629_n4735;
   wire FE_OFN628_n4735;
   wire FE_OFN627_n4735;
   wire FE_OFN626_n4735;
   wire FE_OFN625_n4735;
   wire FE_OFN624_n4735;
   wire FE_OFN623_n4735;
   wire FE_OFN622_n4735;
   wire FE_OFN621_n4735;
   wire FE_OFN620_n4735;
   wire FE_OFN619_n4735;
   wire FE_OFN618_n4735;
   wire FE_OFN617_n4729;
   wire FE_OFN616_n4729;
   wire FE_OFN615_n4729;
   wire FE_OFN614_n4729;
   wire FE_OFN613_n4729;
   wire FE_OFN612_n4729;
   wire FE_OFN611_n4729;
   wire FE_OFN610_n4729;
   wire FE_OFN609_n4729;
   wire FE_OFN608_n4729;
   wire FE_OFN607_n4729;
   wire FE_OFN606_n4729;
   wire FE_OFN605_n4723;
   wire FE_OFN604_n4723;
   wire FE_OFN603_n4723;
   wire FE_OFN602_n4723;
   wire FE_OFN601_n4723;
   wire FE_OFN600_n4723;
   wire FE_OFN599_n4723;
   wire FE_OFN598_n4723;
   wire FE_OFN597_n4723;
   wire FE_OFN596_n4723;
   wire FE_OFN595_n4723;
   wire FE_OFN594_n4723;
   wire FE_OFN593_n4723;
   wire FE_OFN592_n4724;
   wire FE_OFN591_n4724;
   wire FE_OFN590_n4724;
   wire FE_OFN589_n4724;
   wire FE_OFN588_n4724;
   wire FE_OFN587_n4724;
   wire FE_OFN586_n4724;
   wire FE_OFN585_n4724;
   wire FE_OFN584_n4724;
   wire FE_OFN583_n4724;
   wire FE_OFN582_n4724;
   wire FE_OFN581_n4717;
   wire FE_OFN580_n4717;
   wire FE_OFN579_n4717;
   wire FE_OFN578_n4717;
   wire FE_OFN577_n4717;
   wire FE_OFN576_n4717;
   wire FE_OFN575_n4717;
   wire FE_OFN574_n4717;
   wire FE_OFN573_n4717;
   wire FE_OFN572_n4717;
   wire FE_OFN571_n4717;
   wire FE_OFN570_n4717;
   wire FE_OFN569_n4711;
   wire FE_OFN568_n4711;
   wire FE_OFN567_n4711;
   wire FE_OFN566_n4711;
   wire FE_OFN565_n4711;
   wire FE_OFN564_n4711;
   wire FE_OFN563_n4711;
   wire FE_OFN562_n4711;
   wire FE_OFN561_n4711;
   wire FE_OFN560_n4711;
   wire FE_OFN559_n4711;
   wire FE_OFN558_n4711;
   wire FE_OFN557_n4705;
   wire FE_OFN556_n4705;
   wire FE_OFN555_n4705;
   wire FE_OFN554_n4705;
   wire FE_OFN553_n4705;
   wire FE_OFN552_n4705;
   wire FE_OFN551_n4705;
   wire FE_OFN550_n4705;
   wire FE_OFN549_n4705;
   wire FE_OFN548_n4705;
   wire FE_OFN547_n4705;
   wire FE_OFN546_n4705;
   wire FE_OFN545_n4699;
   wire FE_OFN544_n4699;
   wire FE_OFN543_n4699;
   wire FE_OFN542_n4699;
   wire FE_OFN541_n4699;
   wire FE_OFN540_n4699;
   wire FE_OFN539_n4699;
   wire FE_OFN538_n4699;
   wire FE_OFN537_n4699;
   wire FE_OFN536_n4699;
   wire FE_OFN535_n4699;
   wire FE_OFN534_n4699;
   wire FE_OFN533_n4700;
   wire FE_OFN532_n4700;
   wire FE_OFN531_n4700;
   wire FE_OFN530_n4700;
   wire FE_OFN529_n4700;
   wire FE_OFN528_n4700;
   wire FE_OFN527_n4700;
   wire FE_OFN526_n4700;
   wire FE_OFN525_n4700;
   wire FE_OFN524_n4700;
   wire FE_OFN523_n4700;
   wire FE_OFN522_n4693;
   wire FE_OFN521_n4693;
   wire FE_OFN520_n4693;
   wire FE_OFN519_n4693;
   wire FE_OFN518_n4693;
   wire FE_OFN517_n4693;
   wire FE_OFN516_n4693;
   wire FE_OFN515_n4693;
   wire FE_OFN514_n4693;
   wire FE_OFN513_n4693;
   wire FE_OFN512_n4693;
   wire FE_OFN511_n4693;
   wire FE_OFN510_n8055;
   wire FE_OFN509_n8055;
   wire FE_OFN508_n8055;
   wire FE_OFN507_n4681;
   wire FE_OFN506_n4681;
   wire FE_OFN505_n4681;
   wire FE_OFN504_n4681;
   wire FE_OFN503_n4681;
   wire FE_OFN502_n4681;
   wire FE_OFN501_n4681;
   wire FE_OFN500_n4681;
   wire FE_OFN499_n4681;
   wire FE_OFN498_n4681;
   wire FE_OFN497_n4681;
   wire FE_OFN496_n4681;
   wire FE_OFN495_n4682;
   wire FE_OFN494_n4682;
   wire FE_OFN493_n4682;
   wire FE_OFN492_n4682;
   wire FE_OFN491_n4682;
   wire FE_OFN490_n4682;
   wire FE_OFN489_n4682;
   wire FE_OFN488_n4682;
   wire FE_OFN487_n4682;
   wire FE_OFN486_n4682;
   wire FE_OFN485_n4675;
   wire FE_OFN484_n4675;
   wire FE_OFN483_n4675;
   wire FE_OFN482_n4675;
   wire FE_OFN481_n4675;
   wire FE_OFN480_n4675;
   wire FE_OFN479_n4675;
   wire FE_OFN478_n4675;
   wire FE_OFN477_n4675;
   wire FE_OFN476_n4675;
   wire FE_OFN475_n4675;
   wire FE_OFN474_n4675;
   wire FE_OFN473_n4676;
   wire FE_OFN472_n4676;
   wire FE_OFN471_n4676;
   wire FE_OFN470_n4676;
   wire FE_OFN469_n4676;
   wire FE_OFN468_n4676;
   wire FE_OFN467_n4676;
   wire FE_OFN466_n4676;
   wire FE_OFN465_n4676;
   wire FE_OFN464_n4676;
   wire FE_OFN463_n4676;
   wire FE_OFN462_n4688;
   wire FE_OFN461_n4688;
   wire FE_OFN460_n4688;
   wire FE_OFN459_n4688;
   wire FE_OFN458_n4688;
   wire FE_OFN457_n4688;
   wire FE_OFN456_n4688;
   wire FE_OFN455_n4688;
   wire FE_OFN454_n4688;
   wire FE_OFN453_n4688;
   wire FE_OFN452_n4694;
   wire FE_OFN451_n4694;
   wire FE_OFN450_n4694;
   wire FE_OFN449_n4694;
   wire FE_OFN448_n4694;
   wire FE_OFN447_n4694;
   wire FE_OFN446_n4694;
   wire FE_OFN445_n4694;
   wire FE_OFN444_n4694;
   wire FE_OFN443_n4694;
   wire FE_OFN442_n4706;
   wire FE_OFN441_n4706;
   wire FE_OFN440_n4706;
   wire FE_OFN439_n4706;
   wire FE_OFN438_n4706;
   wire FE_OFN437_n4706;
   wire FE_OFN436_n4706;
   wire FE_OFN435_n4706;
   wire FE_OFN434_n4706;
   wire FE_OFN433_n4706;
   wire FE_OFN432_n4712;
   wire FE_OFN431_n4712;
   wire FE_OFN430_n4712;
   wire FE_OFN429_n4712;
   wire FE_OFN428_n4712;
   wire FE_OFN427_n4712;
   wire FE_OFN426_n4712;
   wire FE_OFN425_n4712;
   wire FE_OFN424_n4712;
   wire FE_OFN423_n4712;
   wire FE_OFN422_n3776;
   wire FE_OFN421_n3776;
   wire FE_OFN420_n3776;
   wire FE_OFN419_n3776;
   wire FE_OFN418_n3776;
   wire FE_OFN417_n3776;
   wire FE_OFN416_n3776;
   wire FE_OFN415_n3776;
   wire FE_OFN414_n3776;
   wire FE_OFN413_n3776;
   wire FE_OFN412_n3776;
   wire FE_OFN411_n3777;
   wire FE_OFN410_n3777;
   wire FE_OFN409_n3777;
   wire FE_OFN408_n3777;
   wire FE_OFN407_n3777;
   wire FE_OFN406_n3777;
   wire FE_OFN405_n3777;
   wire FE_OFN404_n3777;
   wire FE_OFN403_n3777;
   wire FE_OFN402_n3777;
   wire FE_OFN401_n3777;
   wire FE_OFN400_n4718;
   wire FE_OFN399_n4718;
   wire FE_OFN398_n4718;
   wire FE_OFN397_n4718;
   wire FE_OFN396_n4718;
   wire FE_OFN395_n4718;
   wire FE_OFN394_n4718;
   wire FE_OFN393_n4718;
   wire FE_OFN392_n4718;
   wire FE_OFN391_n4718;
   wire FE_OFN390_n4718;
   wire FE_OFN389_n4730;
   wire FE_OFN388_n4730;
   wire FE_OFN387_n4730;
   wire FE_OFN386_n4730;
   wire FE_OFN385_n4730;
   wire FE_OFN384_n4730;
   wire FE_OFN383_n4730;
   wire FE_OFN382_n4730;
   wire FE_OFN381_n4730;
   wire FE_OFN380_n4730;
   wire FE_OFN379_n4730;
   wire FE_OFN378_n4736;
   wire FE_OFN377_n4736;
   wire FE_OFN376_n4736;
   wire FE_OFN375_n4736;
   wire FE_OFN374_n4736;
   wire FE_OFN373_n4736;
   wire FE_OFN372_n4736;
   wire FE_OFN371_n4736;
   wire FE_OFN370_n4736;
   wire FE_OFN369_n4736;
   wire FE_OFN368_n4748;
   wire FE_OFN367_n4748;
   wire FE_OFN366_n4748;
   wire FE_OFN365_n4748;
   wire FE_OFN364_n4748;
   wire FE_OFN363_n4748;
   wire FE_OFN362_n4748;
   wire FE_OFN361_n4748;
   wire FE_OFN360_n4748;
   wire FE_OFN359_n4748;
   wire FE_OFN358_n4754;
   wire FE_OFN357_n4754;
   wire FE_OFN356_n4754;
   wire FE_OFN355_n4754;
   wire FE_OFN354_n4754;
   wire FE_OFN353_n4754;
   wire FE_OFN352_n4754;
   wire FE_OFN351_n4754;
   wire FE_OFN350_n4754;
   wire FE_OFN349_n4754;
   wire FE_OFN348_n4760;
   wire FE_OFN347_n4760;
   wire FE_OFN346_n4760;
   wire FE_OFN345_n4760;
   wire FE_OFN344_n4760;
   wire FE_OFN343_n4760;
   wire FE_OFN342_n4760;
   wire FE_OFN341_n4760;
   wire FE_OFN340_n4760;
   wire FE_OFN339_n4760;
   wire FE_OFN338_n4760;
   wire FE_OFN337_n4573;
   wire FE_OFN336_n4573;
   wire FE_OFN335_n4573;
   wire FE_OFN334_n4573;
   wire FE_OFN333_n4573;
   wire FE_OFN332_n4573;
   wire FE_OFN331_n4573;
   wire FE_OFN330_n4573;
   wire FE_OFN329_n4573;
   wire FE_OFN328_n4573;
   wire FE_OFN327_n4573;
   wire FE_OFN326_n8056;
   wire FE_OFN325_n8056;
   wire FE_OFN324_n4561;
   wire FE_OFN323_n4561;
   wire FE_OFN322_n4561;
   wire FE_OFN321_n4561;
   wire FE_OFN320_n4561;
   wire FE_OFN319_n4561;
   wire FE_OFN318_n4561;
   wire FE_OFN317_n4561;
   wire FE_OFN316_n4561;
   wire FE_OFN315_n4561;
   wire FE_OFN314_n4561;
   wire FE_OFN313_n4561;
   wire FE_OFN312_n4555;
   wire FE_OFN311_n4555;
   wire FE_OFN310_n4555;
   wire FE_OFN309_n4555;
   wire FE_OFN308_n4555;
   wire FE_OFN307_n4555;
   wire FE_OFN306_n4555;
   wire FE_OFN305_n4555;
   wire FE_OFN304_n4555;
   wire FE_OFN303_n4555;
   wire FE_OFN302_n4555;
   wire FE_OFN301_n4555;
   wire FE_OFN300_n4556;
   wire FE_OFN299_n4556;
   wire FE_OFN298_n4556;
   wire FE_OFN297_n4556;
   wire FE_OFN296_n4556;
   wire FE_OFN295_n4556;
   wire FE_OFN294_n4556;
   wire FE_OFN293_n4556;
   wire FE_OFN292_n4556;
   wire FE_OFN291_n4556;
   wire FE_OFN290_n4549;
   wire FE_OFN289_n4549;
   wire FE_OFN288_n4549;
   wire FE_OFN287_n4549;
   wire FE_OFN286_n4549;
   wire FE_OFN285_n4549;
   wire FE_OFN284_n4549;
   wire FE_OFN283_n4549;
   wire FE_OFN282_n4549;
   wire FE_OFN281_n4549;
   wire FE_OFN280_n4549;
   wire FE_OFN279_n4549;
   wire FE_OFN278_n4543;
   wire FE_OFN277_n4543;
   wire FE_OFN276_n4543;
   wire FE_OFN275_n4543;
   wire FE_OFN274_n4543;
   wire FE_OFN273_n4543;
   wire FE_OFN272_n4543;
   wire FE_OFN271_n4543;
   wire FE_OFN270_n4543;
   wire FE_OFN269_n4543;
   wire FE_OFN268_n4543;
   wire FE_OFN267_n4543;
   wire FE_OFN266_n4543;
   wire FE_OFN265_n4544;
   wire FE_OFN264_n4544;
   wire FE_OFN263_n4544;
   wire FE_OFN262_n4544;
   wire FE_OFN261_n4544;
   wire FE_OFN260_n4544;
   wire FE_OFN259_n4544;
   wire FE_OFN258_n4544;
   wire FE_OFN257_n4544;
   wire FE_OFN256_n4544;
   wire FE_OFN255_n4537;
   wire FE_OFN254_n4537;
   wire FE_OFN253_n4537;
   wire FE_OFN252_n4537;
   wire FE_OFN251_n4537;
   wire FE_OFN250_n4537;
   wire FE_OFN249_n4537;
   wire FE_OFN248_n4537;
   wire FE_OFN247_n4537;
   wire FE_OFN246_n4537;
   wire FE_OFN245_n4537;
   wire FE_OFN244_n4537;
   wire FE_OFN243_n4531;
   wire FE_OFN242_n4531;
   wire FE_OFN241_n4531;
   wire FE_OFN240_n4531;
   wire FE_OFN239_n4531;
   wire FE_OFN238_n4531;
   wire FE_OFN237_n4531;
   wire FE_OFN236_n4531;
   wire FE_OFN235_n4531;
   wire FE_OFN234_n4531;
   wire FE_OFN233_n4531;
   wire FE_OFN232_n4531;
   wire FE_OFN231_n4525;
   wire FE_OFN230_n4525;
   wire FE_OFN229_n4525;
   wire FE_OFN228_n4525;
   wire FE_OFN227_n4525;
   wire FE_OFN226_n4525;
   wire FE_OFN225_n4525;
   wire FE_OFN224_n4525;
   wire FE_OFN223_n4525;
   wire FE_OFN222_n4525;
   wire FE_OFN221_n4525;
   wire FE_OFN220_n4519;
   wire FE_OFN219_n4519;
   wire FE_OFN218_n4519;
   wire FE_OFN217_n4519;
   wire FE_OFN216_n4519;
   wire FE_OFN215_n4519;
   wire FE_OFN214_n4519;
   wire FE_OFN213_n4519;
   wire FE_OFN212_n4519;
   wire FE_OFN211_n4519;
   wire FE_OFN210_n4519;
   wire FE_OFN209_n4519;
   wire FE_OFN208_n4513;
   wire FE_OFN207_n4513;
   wire FE_OFN206_n4513;
   wire FE_OFN205_n4513;
   wire FE_OFN204_n4513;
   wire FE_OFN203_n4513;
   wire FE_OFN202_n4513;
   wire FE_OFN201_n4513;
   wire FE_OFN200_n4513;
   wire FE_OFN199_n4513;
   wire FE_OFN198_n4513;
   wire FE_OFN197_n4513;
   wire FE_OFN196_n4514;
   wire FE_OFN195_n4514;
   wire FE_OFN194_n4514;
   wire FE_OFN193_n4514;
   wire FE_OFN192_n4514;
   wire FE_OFN191_n4514;
   wire FE_OFN190_n4514;
   wire FE_OFN189_n4514;
   wire FE_OFN188_n4514;
   wire FE_OFN187_n4514;
   wire FE_OFN186_n4507;
   wire FE_OFN185_n4507;
   wire FE_OFN184_n4507;
   wire FE_OFN183_n4507;
   wire FE_OFN182_n4507;
   wire FE_OFN181_n4507;
   wire FE_OFN180_n4507;
   wire FE_OFN179_n4507;
   wire FE_OFN178_n4507;
   wire FE_OFN177_n4507;
   wire FE_OFN176_n4507;
   wire FE_OFN175_n4507;
   wire FE_OFN174_n8054;
   wire FE_OFN173_n8054;
   wire FE_OFN172_n4495;
   wire FE_OFN171_n4495;
   wire FE_OFN170_n4495;
   wire FE_OFN169_n4495;
   wire FE_OFN168_n4495;
   wire FE_OFN167_n4495;
   wire FE_OFN166_n4495;
   wire FE_OFN165_n4495;
   wire FE_OFN164_n4495;
   wire FE_OFN163_n4495;
   wire FE_OFN162_n4495;
   wire FE_OFN161_n4495;
   wire FE_OFN160_n4496;
   wire FE_OFN159_n4496;
   wire FE_OFN158_n4496;
   wire FE_OFN157_n4496;
   wire FE_OFN156_n4496;
   wire FE_OFN155_n4496;
   wire FE_OFN154_n4496;
   wire FE_OFN153_n4496;
   wire FE_OFN152_n4496;
   wire FE_OFN151_n4496;
   wire FE_OFN150_n4489;
   wire FE_OFN149_n4489;
   wire FE_OFN148_n4489;
   wire FE_OFN147_n4489;
   wire FE_OFN146_n4489;
   wire FE_OFN145_n4489;
   wire FE_OFN144_n4489;
   wire FE_OFN143_n4489;
   wire FE_OFN142_n4489;
   wire FE_OFN141_n4489;
   wire FE_OFN140_n4489;
   wire FE_OFN139_n4489;
   wire FE_OFN138_n4490;
   wire FE_OFN137_n4490;
   wire FE_OFN136_n4490;
   wire FE_OFN135_n4490;
   wire FE_OFN134_n4490;
   wire FE_OFN133_n4490;
   wire FE_OFN132_n4490;
   wire FE_OFN131_n4490;
   wire FE_OFN130_n4490;
   wire FE_OFN129_n4490;
   wire FE_OFN128_n4502;
   wire FE_OFN127_n4502;
   wire FE_OFN126_n4502;
   wire FE_OFN125_n4502;
   wire FE_OFN124_n4502;
   wire FE_OFN123_n4502;
   wire FE_OFN122_n4502;
   wire FE_OFN121_n4502;
   wire FE_OFN120_n4502;
   wire FE_OFN119_n4502;
   wire FE_OFN118_n4502;
   wire FE_OFN117_n4502;
   wire FE_OFN116_n4502;
   wire FE_OFN115_n4502;
   wire FE_OFN114_n4508;
   wire FE_OFN113_n4508;
   wire FE_OFN112_n4508;
   wire FE_OFN111_n4508;
   wire FE_OFN110_n4508;
   wire FE_OFN109_n4508;
   wire FE_OFN108_n4508;
   wire FE_OFN107_n4508;
   wire FE_OFN106_n4508;
   wire FE_OFN105_n4508;
   wire FE_OFN104_n4520;
   wire FE_OFN103_n4520;
   wire FE_OFN102_n4520;
   wire FE_OFN101_n4520;
   wire FE_OFN100_n4520;
   wire FE_OFN99_n4520;
   wire FE_OFN98_n4520;
   wire FE_OFN97_n4520;
   wire FE_OFN96_n4520;
   wire FE_OFN95_n4520;
   wire FE_OFN94_n4526;
   wire FE_OFN93_n4526;
   wire FE_OFN92_n4526;
   wire FE_OFN91_n4526;
   wire FE_OFN90_n4526;
   wire FE_OFN89_n4526;
   wire FE_OFN88_n4526;
   wire FE_OFN87_n4526;
   wire FE_OFN86_n4526;
   wire FE_OFN85_n4526;
   wire FE_OFN84_n4526;
   wire FE_OFN83_n3796;
   wire FE_OFN82_n3796;
   wire FE_OFN81_n3796;
   wire FE_OFN80_n3796;
   wire FE_OFN79_n3796;
   wire FE_OFN78_n3796;
   wire FE_OFN77_n3796;
   wire FE_OFN76_n3796;
   wire FE_OFN75_n3796;
   wire FE_OFN74_n3796;
   wire FE_OFN73_n3796;
   wire FE_OFN72_n3797;
   wire FE_OFN71_n3797;
   wire FE_OFN70_n3797;
   wire FE_OFN69_n3797;
   wire FE_OFN68_n3797;
   wire FE_OFN67_n3797;
   wire FE_OFN66_n3797;
   wire FE_OFN65_n3797;
   wire FE_OFN64_n3797;
   wire FE_OFN63_n3797;
   wire FE_OFN62_n4532;
   wire FE_OFN61_n4532;
   wire FE_OFN60_n4532;
   wire FE_OFN59_n4532;
   wire FE_OFN58_n4532;
   wire FE_OFN57_n4532;
   wire FE_OFN56_n4532;
   wire FE_OFN55_n4532;
   wire FE_OFN54_n4532;
   wire FE_OFN53_n4532;
   wire FE_OFN52_n4538;
   wire FE_OFN51_n4538;
   wire FE_OFN50_n4538;
   wire FE_OFN49_n4538;
   wire FE_OFN48_n4538;
   wire FE_OFN47_n4538;
   wire FE_OFN46_n4538;
   wire FE_OFN45_n4538;
   wire FE_OFN44_n4538;
   wire FE_OFN43_n4538;
   wire FE_OFN42_n4550;
   wire FE_OFN41_n4550;
   wire FE_OFN40_n4550;
   wire FE_OFN39_n4550;
   wire FE_OFN38_n4550;
   wire FE_OFN37_n4550;
   wire FE_OFN36_n4550;
   wire FE_OFN35_n4550;
   wire FE_OFN34_n4550;
   wire FE_OFN33_n4550;
   wire FE_OFN32_n4562;
   wire FE_OFN31_n4562;
   wire FE_OFN30_n4562;
   wire FE_OFN29_n4562;
   wire FE_OFN28_n4562;
   wire FE_OFN27_n4562;
   wire FE_OFN26_n4562;
   wire FE_OFN25_n4562;
   wire FE_OFN24_n4562;
   wire FE_OFN23_n4562;
   wire FE_OFN22_n4562;
   wire FE_OFN21_n4568;
   wire FE_OFN20_n4568;
   wire FE_OFN19_n4568;
   wire FE_OFN18_n4568;
   wire FE_OFN17_n4568;
   wire FE_OFN16_n4568;
   wire FE_OFN15_n4568;
   wire FE_OFN14_n4568;
   wire FE_OFN13_n4568;
   wire FE_OFN12_n4568;
   wire FE_OFN11_n4568;
   wire FE_OFN10_n4568;
   wire FE_OFN9_n4574;
   wire FE_OFN8_n4574;
   wire FE_OFN7_n4574;
   wire FE_OFN6_n4574;
   wire FE_OFN5_n4574;
   wire FE_OFN4_n4574;
   wire FE_OFN3_n4574;
   wire FE_OFN2_n4574;
   wire FE_OFN1_n4574;
   wire FE_OFN0_n4574;
   wire FE_MDBN14_;
   wire FE_MDBN13_;
   wire FE_MDBN12_;
   wire FE_MDBN11_;
   wire FE_MDBN10_;
   wire FE_MDBN9_;
   wire FE_MDBN8_;
   wire FE_MDBN7_;
   wire FE_MDBN6_;
   wire FE_MDBN5_;
   wire FE_MDBN4_;
   wire FE_MDBN3_;
   wire FE_MDBN2_;
   wire FE_MDBN1_;
   wire FE_MDBN0_;
   wire n9614;
   wire n9615;
   wire acc_done;
   wire acc_bypass;
   wire from_fft_empty;
   wire from_fir_empty;
   wire iir_enable;
   wire \fifo_to_fft/hang[14] ;
   wire \fifo_to_fft/hang[13] ;
   wire \fifo_to_fft/hang[12] ;
   wire \fifo_to_fft/hang[11] ;
   wire \fifo_to_fft/hang[10] ;
   wire \fifo_to_fft/hang[9] ;
   wire \fifo_to_fft/hang[8] ;
   wire \fifo_to_fft/hang[7] ;
   wire \fifo_to_fft/hang[6] ;
   wire \fifo_to_fft/hang[5] ;
   wire \fifo_to_fft/hang[4] ;
   wire \fifo_to_fft/hang[3] ;
   wire \fifo_to_fft/hang[2] ;
   wire \fifo_to_fft/hang[1] ;
   wire \fifo_to_fft/hang[0] ;
   wire \fifo_to_fft/hold[15] ;
   wire \fifo_to_fft/hold[14] ;
   wire \fifo_to_fft/hold[13] ;
   wire \fifo_to_fft/hold[12] ;
   wire \fifo_to_fft/hold[11] ;
   wire \fifo_to_fft/hold[10] ;
   wire \fifo_to_fft/hold[9] ;
   wire \fifo_to_fft/hold[8] ;
   wire \fifo_to_fft/hold[7] ;
   wire \fifo_to_fft/hold[6] ;
   wire \fifo_to_fft/hold[5] ;
   wire \fifo_to_fft/hold[4] ;
   wire \fifo_to_fft/hold[3] ;
   wire \fifo_to_fft/hold[2] ;
   wire \fifo_to_fft/hold[1] ;
   wire \fifo_to_fft/hold[0] ;
   wire \fifo_to_fft/tok_xnor_put ;
   wire \fifo_from_fft/hang[14] ;
   wire \fifo_from_fft/hang[13] ;
   wire \fifo_from_fft/hang[12] ;
   wire \fifo_from_fft/hang[11] ;
   wire \fifo_from_fft/hang[10] ;
   wire \fifo_from_fft/hang[9] ;
   wire \fifo_from_fft/hang[8] ;
   wire \fifo_from_fft/hang[7] ;
   wire \fifo_from_fft/hang[6] ;
   wire \fifo_from_fft/hang[5] ;
   wire \fifo_from_fft/hang[4] ;
   wire \fifo_from_fft/hang[3] ;
   wire \fifo_from_fft/hang[2] ;
   wire \fifo_from_fft/hang[1] ;
   wire \fifo_from_fft/hang[0] ;
   wire \fifo_from_fft/hold[15] ;
   wire \fifo_from_fft/hold[14] ;
   wire \fifo_from_fft/hold[13] ;
   wire \fifo_from_fft/hold[12] ;
   wire \fifo_from_fft/hold[11] ;
   wire \fifo_from_fft/hold[10] ;
   wire \fifo_from_fft/hold[9] ;
   wire \fifo_from_fft/hold[8] ;
   wire \fifo_from_fft/hold[7] ;
   wire \fifo_from_fft/hold[6] ;
   wire \fifo_from_fft/hold[5] ;
   wire \fifo_from_fft/hold[4] ;
   wire \fifo_from_fft/hold[3] ;
   wire \fifo_from_fft/hold[2] ;
   wire \fifo_from_fft/hold[1] ;
   wire \fifo_from_fft/hold[0] ;
   wire \fifo_from_fft/tok_xnor_put ;
   wire \fifo_to_fir/hang[14] ;
   wire \fifo_to_fir/hang[13] ;
   wire \fifo_to_fir/hang[12] ;
   wire \fifo_to_fir/hang[11] ;
   wire \fifo_to_fir/hang[10] ;
   wire \fifo_to_fir/hang[9] ;
   wire \fifo_to_fir/hang[8] ;
   wire \fifo_to_fir/hang[7] ;
   wire \fifo_to_fir/hang[6] ;
   wire \fifo_to_fir/hang[5] ;
   wire \fifo_to_fir/hang[4] ;
   wire \fifo_to_fir/hang[3] ;
   wire \fifo_to_fir/hang[2] ;
   wire \fifo_to_fir/hang[1] ;
   wire \fifo_to_fir/hang[0] ;
   wire \fifo_to_fir/hold[15] ;
   wire \fifo_to_fir/hold[14] ;
   wire \fifo_to_fir/hold[13] ;
   wire \fifo_to_fir/hold[12] ;
   wire \fifo_to_fir/hold[11] ;
   wire \fifo_to_fir/hold[10] ;
   wire \fifo_to_fir/hold[9] ;
   wire \fifo_to_fir/hold[8] ;
   wire \fifo_to_fir/hold[7] ;
   wire \fifo_to_fir/hold[6] ;
   wire \fifo_to_fir/hold[5] ;
   wire \fifo_to_fir/hold[4] ;
   wire \fifo_to_fir/hold[3] ;
   wire \fifo_to_fir/hold[2] ;
   wire \fifo_to_fir/hold[1] ;
   wire \fifo_to_fir/hold[0] ;
   wire \fifo_to_fir/tok_xnor_put ;
   wire \fifo_from_fir/hang[14] ;
   wire \fifo_from_fir/hang[13] ;
   wire \fifo_from_fir/hang[12] ;
   wire \fifo_from_fir/hang[11] ;
   wire \fifo_from_fir/hang[10] ;
   wire \fifo_from_fir/hang[9] ;
   wire \fifo_from_fir/hang[8] ;
   wire \fifo_from_fir/hang[7] ;
   wire \fifo_from_fir/hang[6] ;
   wire \fifo_from_fir/hang[5] ;
   wire \fifo_from_fir/hang[4] ;
   wire \fifo_from_fir/hang[3] ;
   wire \fifo_from_fir/hang[2] ;
   wire \fifo_from_fir/hang[1] ;
   wire \fifo_from_fir/hang[0] ;
   wire \fifo_from_fir/hold[15] ;
   wire \fifo_from_fir/hold[14] ;
   wire \fifo_from_fir/hold[13] ;
   wire \fifo_from_fir/hold[12] ;
   wire \fifo_from_fir/hold[11] ;
   wire \fifo_from_fir/hold[10] ;
   wire \fifo_from_fir/hold[9] ;
   wire \fifo_from_fir/hold[8] ;
   wire \fifo_from_fir/hold[7] ;
   wire \fifo_from_fir/hold[6] ;
   wire \fifo_from_fir/hold[5] ;
   wire \fifo_from_fir/hold[4] ;
   wire \fifo_from_fir/hold[3] ;
   wire \fifo_from_fir/hold[2] ;
   wire \fifo_from_fir/hold[1] ;
   wire \fifo_from_fir/hold[0] ;
   wire \fifo_from_fir/tok_xnor_put ;
   wire \router/ram_write_enable_reg ;
   wire \router/ram_read_enable_reg ;
   wire \router/iir_get_req_reg ;
   wire \router/fir_get_req_reg ;
   wire \router/fir_put_req_reg ;
   wire \router/fft_get_req_reg ;
   wire \router/fft_put_req_reg ;
   wire \router/iir_write_done ;
   wire \router/fir_write_done ;
   wire \router/fir_read_done ;
   wire \router/fft_write_done ;
   wire \router/fft_read_done ;
   wire \router/data_from_iir ;
   wire \router/data_from_fir ;
   wire \router/data_to_fir ;
   wire \router/data_from_fft ;
   wire \router/data_to_fft ;
   wire \mips/mips/accfullinstruction[31] ;
   wire \mips/mips/accfullinstruction[30] ;
   wire \mips/mips/accfullinstruction[29] ;
   wire \mips/mips/accfullinstruction[28] ;
   wire \mips/mips/accfullinstruction[27] ;
   wire \mips/mips/accfullinstruction[26] ;
   wire \mips/mips/accfullinstruction[25] ;
   wire \mips/mips/accfullinstruction[24] ;
   wire \mips/mips/accfullinstruction[23] ;
   wire \mips/mips/accfullinstruction[22] ;
   wire \mips/mips/accfullinstruction[21] ;
   wire \mips/mips/accfullinstruction[20] ;
   wire \mips/mips/accfullinstruction[19] ;
   wire \mips/mips/accfullinstruction[18] ;
   wire \mips/mips/accfullinstruction[17] ;
   wire \mips/mips/accfullinstruction[16] ;
   wire \mips/mips/accfullinstruction[15] ;
   wire \mips/mips/accfullinstruction[14] ;
   wire \mips/mips/accfullinstruction[13] ;
   wire \mips/mips/accfullinstruction[12] ;
   wire \mips/mips/accfullinstruction[11] ;
   wire \mips/mips/accfullinstruction[10] ;
   wire \mips/mips/accfullinstruction[9] ;
   wire \mips/mips/accfullinstruction[8] ;
   wire \mips/mips/accfullinstruction[7] ;
   wire \mips/mips/accfullinstruction[6] ;
   wire \mips/mips/accfullinstruction[5] ;
   wire \mips/mips/accfullinstruction[4] ;
   wire \mips/mips/accfullinstruction[3] ;
   wire \mips/mips/accfullinstruction[2] ;
   wire \mips/mips/accfullinstruction[1] ;
   wire \mips/mips/accfullinstruction[0] ;
   wire \mips/mips/accbypass ;
   wire \fifo_to_fft/fifo_cell0/N7 ;
   wire \fifo_to_fft/fifo_cell0/control_signal ;
   wire \fifo_to_fft/fifo_cell15/N7 ;
   wire \fifo_to_fft/fifo_cell15/control_signal ;
   wire \fifo_to_fft/empty_det/N4 ;
   wire \fifo_from_fft/fifo_cell0/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell0/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell1/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell2/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell3/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell4/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell5/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell6/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell7/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell8/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell9/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell10/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell11/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell12/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell13/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell14/sr_out[0] ;
   wire \fifo_from_fft/fifo_cell15/N7 ;
   wire \fifo_from_fft/fifo_cell15/sr_out[31] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[30] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[29] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[28] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[27] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[26] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[25] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[24] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[23] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[22] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[21] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[20] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[19] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[18] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[17] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[16] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[15] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[14] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[13] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[12] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[11] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[10] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[9] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[8] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[7] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[6] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[5] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[4] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[3] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[2] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[1] ;
   wire \fifo_from_fft/fifo_cell15/sr_out[0] ;
   wire \fifo_from_fft/empty_det/N4 ;
   wire \fifo_to_fir/fifo_cell0/N7 ;
   wire \fifo_to_fir/fifo_cell0/control_signal ;
   wire \fifo_to_fir/fifo_cell15/N7 ;
   wire \fifo_to_fir/fifo_cell15/control_signal ;
   wire \fifo_to_fir/empty_det/N4 ;
   wire \fifo_from_fir/fifo_cell0/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell0/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell1/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell2/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell3/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell4/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell5/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell6/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell7/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell8/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell9/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell10/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell11/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell12/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell13/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell14/sr_out[0] ;
   wire \fifo_from_fir/fifo_cell15/N7 ;
   wire \fifo_from_fir/fifo_cell15/sr_out[31] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[30] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[29] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[28] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[27] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[26] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[25] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[24] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[23] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[22] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[21] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[20] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[19] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[18] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[17] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[16] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[15] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[14] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[13] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[12] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[11] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[10] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[9] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[8] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[7] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[6] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[5] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[4] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[3] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[2] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[1] ;
   wire \fifo_from_fir/fifo_cell15/sr_out[0] ;
   wire \fifo_from_fir/empty_det/N4 ;
   wire \router/pla_top/N60 ;
   wire \router/pla_top/instruction_valid ;
   wire \router/addr_calc/N191 ;
   wire \router/addr_calc/N99 ;
   wire \router/addr_calc/N95 ;
   wire \router/addr_calc/N63 ;
   wire \router/addr_calc/N9 ;
   wire \router/data_cntl/data_in[31] ;
   wire \router/data_cntl/data_in[30] ;
   wire \router/data_cntl/data_in[29] ;
   wire \router/data_cntl/data_in[28] ;
   wire \router/data_cntl/data_in[27] ;
   wire \router/data_cntl/data_in[26] ;
   wire \router/data_cntl/data_in[25] ;
   wire \router/data_cntl/data_in[24] ;
   wire \router/data_cntl/data_in[23] ;
   wire \router/data_cntl/data_in[22] ;
   wire \router/data_cntl/data_in[21] ;
   wire \router/data_cntl/data_in[20] ;
   wire \router/data_cntl/data_in[19] ;
   wire \router/data_cntl/data_in[18] ;
   wire \router/data_cntl/data_in[17] ;
   wire \router/data_cntl/data_in[16] ;
   wire \router/data_cntl/data_in[15] ;
   wire \router/data_cntl/data_in[14] ;
   wire \router/data_cntl/data_in[13] ;
   wire \router/data_cntl/data_in[12] ;
   wire \router/data_cntl/data_in[11] ;
   wire \router/data_cntl/data_in[10] ;
   wire \router/data_cntl/data_in[9] ;
   wire \router/data_cntl/data_in[8] ;
   wire \router/data_cntl/data_in[7] ;
   wire \router/data_cntl/data_in[6] ;
   wire \router/data_cntl/data_in[5] ;
   wire \router/data_cntl/data_in[4] ;
   wire \router/data_cntl/data_in[3] ;
   wire \router/data_cntl/data_in[2] ;
   wire \router/data_cntl/data_in[1] ;
   wire \router/data_cntl/data_in[0] ;
   wire \router/data_cntl/N151 ;
   wire \router/data_cntl/N142 ;
   wire \router/data_cntl/N139 ;
   wire \router/data_cntl/N138 ;
   wire \router/data_cntl/N137 ;
   wire \router/data_cntl/N135 ;
   wire \router/data_cntl/N134 ;
   wire \router/data_cntl/N133 ;
   wire \router/data_cntl/fir_full_flag ;
   wire \router/data_cntl/fft_full_flag ;
   wire \mips/mips/a/N50 ;
   wire \mips/mips/a/N49 ;
   wire \mips/mips/a/countflag ;
   wire \mips/mips/a/count[0] ;
   wire \fifo_to_fft/fifo_cell0/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell0/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell0/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell0/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell0/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell0/reg_ptok/N22 ;
   wire \fifo_to_fft/fifo_cell0/reg_ptok/out_valid_get ;
   wire \fifo_to_fft/fifo_cell0/reg_ptok/out_valid_put ;
   wire \fifo_to_fft/fifo_cell0/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell1/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell1/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell1/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell1/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell1/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell1/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell2/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell2/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell2/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell2/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell2/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell2/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell3/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell3/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell3/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell3/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell3/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell3/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell4/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell4/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell4/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell4/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell4/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell4/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell5/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell5/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell5/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell5/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell5/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell5/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell6/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell6/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell6/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell6/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell6/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell6/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell7/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell7/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell7/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell7/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell7/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell7/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell8/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell8/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell8/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell8/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell8/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell8/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell9/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell9/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell9/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell9/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell9/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell9/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell10/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell10/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell10/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell10/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell10/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell10/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell11/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell11/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell11/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell11/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell11/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell11/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell12/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell12/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell12/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell12/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell12/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell12/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell13/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell13/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell13/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell13/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell13/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell13/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell14/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell14/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell14/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell14/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell14/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell14/reg_gtok/token ;
   wire \fifo_to_fft/fifo_cell15/controller/f_i_get ;
   wire \fifo_to_fft/fifo_cell15/controller/valid_read ;
   wire \fifo_to_fft/fifo_cell15/controller/f_i_put ;
   wire \fifo_to_fft/fifo_cell15/controller/write_enable ;
   wire \fifo_to_fft/fifo_cell15/data_out/N35 ;
   wire \fifo_to_fft/fifo_cell15/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell0/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell0/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell0/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell0/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell0/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell0/reg_ptok/out_valid_get ;
   wire \fifo_from_fft/fifo_cell0/reg_ptok/out_valid_put ;
   wire \fifo_from_fft/fifo_cell0/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell1/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell1/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell1/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell1/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell1/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell1/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell1/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell2/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell2/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell2/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell2/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell2/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell2/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell2/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell3/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell3/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell3/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell3/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell3/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell3/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell3/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell4/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell4/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell4/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell4/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell4/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell4/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell4/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell5/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell5/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell5/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell5/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell5/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell5/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell5/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell6/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell6/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell6/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell6/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell6/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell6/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell6/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell7/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell7/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell7/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell7/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell7/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell7/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell7/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell8/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell8/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell8/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell8/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell8/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell8/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell8/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell9/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell9/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell9/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell9/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell9/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell9/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell9/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell10/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell10/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell10/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell10/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell10/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell10/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell10/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell11/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell11/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell11/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell11/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell11/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell11/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell11/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell12/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell12/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell12/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell12/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell12/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell12/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell12/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell13/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell13/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell13/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell13/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell13/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell13/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell13/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell14/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell14/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell14/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell14/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell14/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell14/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell14/reg_gtok/token ;
   wire \fifo_from_fft/fifo_cell15/controller/f_i_get ;
   wire \fifo_from_fft/fifo_cell15/controller/valid_read ;
   wire \fifo_from_fft/fifo_cell15/controller/f_i_put ;
   wire \fifo_from_fft/fifo_cell15/controller/write_enable ;
   wire \fifo_from_fft/fifo_cell15/data_out/N35 ;
   wire \fifo_from_fft/fifo_cell15/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell15/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell0/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell0/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell0/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell0/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell0/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell0/reg_ptok/N22 ;
   wire \fifo_to_fir/fifo_cell0/reg_ptok/out_valid_get ;
   wire \fifo_to_fir/fifo_cell0/reg_ptok/out_valid_put ;
   wire \fifo_to_fir/fifo_cell0/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell1/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell1/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell1/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell1/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell1/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell1/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell2/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell2/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell2/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell2/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell2/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell2/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell3/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell3/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell3/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell3/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell3/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell3/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell4/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell4/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell4/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell4/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell4/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell4/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell5/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell5/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell5/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell5/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell5/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell5/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell6/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell6/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell6/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell6/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell6/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell6/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell7/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell7/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell7/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell7/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell7/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell7/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell8/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell8/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell8/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell8/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell8/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell8/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell9/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell9/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell9/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell9/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell9/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell9/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell10/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell10/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell10/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell10/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell10/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell10/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell11/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell11/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell11/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell11/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell11/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell11/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell12/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell12/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell12/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell12/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell12/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell12/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell13/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell13/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell13/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell13/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell13/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell13/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell14/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell14/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell14/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell14/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell14/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell14/reg_gtok/token ;
   wire \fifo_to_fir/fifo_cell15/controller/f_i_get ;
   wire \fifo_to_fir/fifo_cell15/controller/valid_read ;
   wire \fifo_to_fir/fifo_cell15/controller/f_i_put ;
   wire \fifo_to_fir/fifo_cell15/controller/write_enable ;
   wire \fifo_to_fir/fifo_cell15/data_out/N35 ;
   wire \fifo_to_fir/fifo_cell15/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell0/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell0/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell0/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell0/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell0/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell0/reg_ptok/out_valid_get ;
   wire \fifo_from_fir/fifo_cell0/reg_ptok/out_valid_put ;
   wire \fifo_from_fir/fifo_cell0/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell1/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell1/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell1/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell1/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell1/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell1/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell1/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell2/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell2/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell2/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell2/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell2/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell2/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell2/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell3/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell3/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell3/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell3/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell3/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell3/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell3/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell4/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell4/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell4/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell4/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell4/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell4/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell4/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell5/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell5/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell5/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell5/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell5/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell5/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell5/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell6/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell6/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell6/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell6/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell6/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell6/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell6/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell7/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell7/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell7/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell7/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell7/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell7/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell7/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell8/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell8/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell8/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell8/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell8/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell8/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell8/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell9/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell9/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell9/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell9/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell9/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell9/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell9/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell10/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell10/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell10/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell10/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell10/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell10/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell10/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell11/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell11/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell11/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell11/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell11/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell11/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell11/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell12/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell12/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell12/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell12/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell12/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell12/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell12/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell13/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell13/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell13/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell13/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell13/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell13/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell13/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell14/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell14/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell14/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell14/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell14/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell14/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell14/reg_gtok/token ;
   wire \fifo_from_fir/fifo_cell15/controller/f_i_get ;
   wire \fifo_from_fir/fifo_cell15/controller/valid_read ;
   wire \fifo_from_fir/fifo_cell15/controller/f_i_put ;
   wire \fifo_from_fir/fifo_cell15/controller/write_enable ;
   wire \fifo_from_fir/fifo_cell15/data_out/N35 ;
   wire \fifo_from_fir/fifo_cell15/data_out/N9 ;
   wire \fifo_from_fir/fifo_cell15/reg_gtok/token ;
   wire \router/addr_calc/fft_read_calc/count[30] ;
   wire \router/addr_calc/fft_read_calc/count[27] ;
   wire \router/addr_calc/fft_read_calc/count[23] ;
   wire \router/addr_calc/fft_read_calc/count[19] ;
   wire \router/addr_calc/fft_read_calc/count[16] ;
   wire \router/addr_calc/fft_read_calc/count[9] ;
   wire \router/addr_calc/fft_read_calc/count[5] ;
   wire \router/addr_calc/fft_read_calc/count[0] ;
   wire \router/addr_calc/fft_write_calc/count[31] ;
   wire \router/addr_calc/fft_write_calc/count[29] ;
   wire \router/addr_calc/fft_write_calc/count[27] ;
   wire \router/addr_calc/fft_write_calc/count[23] ;
   wire \router/addr_calc/fft_write_calc/count[19] ;
   wire \router/addr_calc/fft_write_calc/count[15] ;
   wire \router/addr_calc/fft_write_calc/count[9] ;
   wire \router/addr_calc/fft_write_calc/count[0] ;
   wire \router/addr_calc/fir_read_calc/count[30] ;
   wire \router/addr_calc/fir_read_calc/count[27] ;
   wire \router/addr_calc/fir_read_calc/count[23] ;
   wire \router/addr_calc/fir_read_calc/count[19] ;
   wire \router/addr_calc/fir_read_calc/count[15] ;
   wire \router/addr_calc/fir_read_calc/count[9] ;
   wire \router/addr_calc/fir_read_calc/count[5] ;
   wire \router/addr_calc/fir_read_calc/count[0] ;
   wire \router/addr_calc/fir_write_calc/count[30] ;
   wire \router/addr_calc/fir_write_calc/count[27] ;
   wire \router/addr_calc/fir_write_calc/count[23] ;
   wire \router/addr_calc/fir_write_calc/count[19] ;
   wire \router/addr_calc/fir_write_calc/count[16] ;
   wire \router/addr_calc/fir_write_calc/count[9] ;
   wire \router/addr_calc/fir_write_calc/count[5] ;
   wire \router/addr_calc/fir_write_calc/count[0] ;
   wire \router/addr_calc/iir_read_calc/count[31] ;
   wire \router/addr_calc/iir_read_calc/count[30] ;
   wire \router/addr_calc/iir_read_calc/count[29] ;
   wire \router/addr_calc/iir_read_calc/count[28] ;
   wire \router/addr_calc/iir_read_calc/count[27] ;
   wire \router/addr_calc/iir_read_calc/count[26] ;
   wire \router/addr_calc/iir_read_calc/count[25] ;
   wire \router/addr_calc/iir_read_calc/count[24] ;
   wire \router/addr_calc/iir_read_calc/count[23] ;
   wire \router/addr_calc/iir_read_calc/count[22] ;
   wire \router/addr_calc/iir_read_calc/count[21] ;
   wire \router/addr_calc/iir_read_calc/count[20] ;
   wire \router/addr_calc/iir_read_calc/count[19] ;
   wire \router/addr_calc/iir_read_calc/count[18] ;
   wire \router/addr_calc/iir_read_calc/count[17] ;
   wire \router/addr_calc/iir_read_calc/count[16] ;
   wire \router/addr_calc/iir_read_calc/count[15] ;
   wire \router/addr_calc/iir_read_calc/count[14] ;
   wire \router/addr_calc/iir_read_calc/count[13] ;
   wire \router/addr_calc/iir_read_calc/count[12] ;
   wire \router/addr_calc/iir_read_calc/count[11] ;
   wire \router/addr_calc/iir_read_calc/count[10] ;
   wire \router/addr_calc/iir_read_calc/count[9] ;
   wire \router/addr_calc/iir_read_calc/count[8] ;
   wire \router/addr_calc/iir_read_calc/count[7] ;
   wire \router/addr_calc/iir_read_calc/count[6] ;
   wire \router/addr_calc/iir_read_calc/count[5] ;
   wire \router/addr_calc/iir_read_calc/count[4] ;
   wire \router/addr_calc/iir_read_calc/count[3] ;
   wire \router/addr_calc/iir_read_calc/count[2] ;
   wire \router/addr_calc/iir_read_calc/count[1] ;
   wire \router/addr_calc/iir_read_calc/count[0] ;
   wire \router/addr_calc/iir_write_calc/count[30] ;
   wire \router/addr_calc/iir_write_calc/count[27] ;
   wire \router/addr_calc/iir_write_calc/count[23] ;
   wire \router/addr_calc/iir_write_calc/count[19] ;
   wire \router/addr_calc/iir_write_calc/count[16] ;
   wire \router/addr_calc/iir_write_calc/count[9] ;
   wire \router/addr_calc/iir_write_calc/count[5] ;
   wire \router/addr_calc/iir_write_calc/count[0] ;
   wire \router/addr_calc/fft_read_calc/counter/N209 ;
   wire \router/addr_calc/fft_read_calc/counter/N208 ;
   wire \router/addr_calc/fft_read_calc/counter/N207 ;
   wire \router/addr_calc/fft_read_calc/counter/N206 ;
   wire \router/addr_calc/fft_read_calc/counter/N205 ;
   wire \router/addr_calc/fft_read_calc/counter/N204 ;
   wire \router/addr_calc/fft_read_calc/counter/N203 ;
   wire \router/addr_calc/fft_read_calc/counter/N202 ;
   wire \router/addr_calc/fft_read_calc/counter/N201 ;
   wire \router/addr_calc/fft_read_calc/counter/N200 ;
   wire \router/addr_calc/fft_read_calc/counter/N199 ;
   wire \router/addr_calc/fft_read_calc/counter/N198 ;
   wire \router/addr_calc/fft_read_calc/counter/N197 ;
   wire \router/addr_calc/fft_read_calc/counter/N196 ;
   wire \router/addr_calc/fft_read_calc/counter/N195 ;
   wire \router/addr_calc/fft_read_calc/counter/N194 ;
   wire \router/addr_calc/fft_read_calc/counter/N193 ;
   wire \router/addr_calc/fft_read_calc/counter/N192 ;
   wire \router/addr_calc/fft_read_calc/counter/N191 ;
   wire \router/addr_calc/fft_read_calc/counter/N190 ;
   wire \router/addr_calc/fft_read_calc/counter/N189 ;
   wire \router/addr_calc/fft_read_calc/counter/N188 ;
   wire \router/addr_calc/fft_read_calc/counter/N187 ;
   wire \router/addr_calc/fft_read_calc/counter/N186 ;
   wire \router/addr_calc/fft_read_calc/counter/N185 ;
   wire \router/addr_calc/fft_read_calc/counter/N184 ;
   wire \router/addr_calc/fft_read_calc/counter/N183 ;
   wire \router/addr_calc/fft_read_calc/counter/N182 ;
   wire \router/addr_calc/fft_read_calc/counter/N181 ;
   wire \router/addr_calc/fft_read_calc/counter/N180 ;
   wire \router/addr_calc/fft_read_calc/counter/N179 ;
   wire \router/addr_calc/fft_read_calc/counter/N178 ;
   wire \router/addr_calc/fft_read_calc/counter/N77 ;
   wire \router/addr_calc/fft_read_calc/counter/N76 ;
   wire \router/addr_calc/fft_read_calc/counter/N75 ;
   wire \router/addr_calc/fft_read_calc/counter/N74 ;
   wire \router/addr_calc/fft_read_calc/counter/N73 ;
   wire \router/addr_calc/fft_read_calc/counter/N72 ;
   wire \router/addr_calc/fft_read_calc/counter/N71 ;
   wire \router/addr_calc/fft_read_calc/counter/N70 ;
   wire \router/addr_calc/fft_read_calc/counter/N69 ;
   wire \router/addr_calc/fft_read_calc/counter/N68 ;
   wire \router/addr_calc/fft_read_calc/counter/N67 ;
   wire \router/addr_calc/fft_read_calc/counter/N66 ;
   wire \router/addr_calc/fft_read_calc/counter/N65 ;
   wire \router/addr_calc/fft_read_calc/counter/N64 ;
   wire \router/addr_calc/fft_read_calc/counter/N63 ;
   wire \router/addr_calc/fft_read_calc/counter/N62 ;
   wire \router/addr_calc/fft_read_calc/counter/N61 ;
   wire \router/addr_calc/fft_read_calc/counter/N60 ;
   wire \router/addr_calc/fft_read_calc/counter/N59 ;
   wire \router/addr_calc/fft_read_calc/counter/N58 ;
   wire \router/addr_calc/fft_read_calc/counter/N57 ;
   wire \router/addr_calc/fft_read_calc/counter/N56 ;
   wire \router/addr_calc/fft_read_calc/counter/N55 ;
   wire \router/addr_calc/fft_read_calc/counter/N54 ;
   wire \router/addr_calc/fft_read_calc/counter/N53 ;
   wire \router/addr_calc/fft_read_calc/counter/N52 ;
   wire \router/addr_calc/fft_read_calc/counter/N51 ;
   wire \router/addr_calc/fft_read_calc/counter/N50 ;
   wire \router/addr_calc/fft_read_calc/counter/N49 ;
   wire \router/addr_calc/fft_read_calc/counter/N48 ;
   wire \router/addr_calc/fft_read_calc/counter/N47 ;
   wire \router/addr_calc/fft_read_calc/counter/N40 ;
   wire \router/addr_calc/fft_read_calc/counter/hold ;
   wire \router/addr_calc/fft_write_calc/counter/N209 ;
   wire \router/addr_calc/fft_write_calc/counter/N208 ;
   wire \router/addr_calc/fft_write_calc/counter/N207 ;
   wire \router/addr_calc/fft_write_calc/counter/N206 ;
   wire \router/addr_calc/fft_write_calc/counter/N205 ;
   wire \router/addr_calc/fft_write_calc/counter/N204 ;
   wire \router/addr_calc/fft_write_calc/counter/N203 ;
   wire \router/addr_calc/fft_write_calc/counter/N202 ;
   wire \router/addr_calc/fft_write_calc/counter/N201 ;
   wire \router/addr_calc/fft_write_calc/counter/N200 ;
   wire \router/addr_calc/fft_write_calc/counter/N199 ;
   wire \router/addr_calc/fft_write_calc/counter/N198 ;
   wire \router/addr_calc/fft_write_calc/counter/N197 ;
   wire \router/addr_calc/fft_write_calc/counter/N196 ;
   wire \router/addr_calc/fft_write_calc/counter/N195 ;
   wire \router/addr_calc/fft_write_calc/counter/N194 ;
   wire \router/addr_calc/fft_write_calc/counter/N193 ;
   wire \router/addr_calc/fft_write_calc/counter/N192 ;
   wire \router/addr_calc/fft_write_calc/counter/N191 ;
   wire \router/addr_calc/fft_write_calc/counter/N190 ;
   wire \router/addr_calc/fft_write_calc/counter/N189 ;
   wire \router/addr_calc/fft_write_calc/counter/N188 ;
   wire \router/addr_calc/fft_write_calc/counter/N187 ;
   wire \router/addr_calc/fft_write_calc/counter/N186 ;
   wire \router/addr_calc/fft_write_calc/counter/N185 ;
   wire \router/addr_calc/fft_write_calc/counter/N184 ;
   wire \router/addr_calc/fft_write_calc/counter/N183 ;
   wire \router/addr_calc/fft_write_calc/counter/N182 ;
   wire \router/addr_calc/fft_write_calc/counter/N181 ;
   wire \router/addr_calc/fft_write_calc/counter/N180 ;
   wire \router/addr_calc/fft_write_calc/counter/N179 ;
   wire \router/addr_calc/fft_write_calc/counter/N178 ;
   wire \router/addr_calc/fft_write_calc/counter/N77 ;
   wire \router/addr_calc/fft_write_calc/counter/N76 ;
   wire \router/addr_calc/fft_write_calc/counter/N75 ;
   wire \router/addr_calc/fft_write_calc/counter/N74 ;
   wire \router/addr_calc/fft_write_calc/counter/N73 ;
   wire \router/addr_calc/fft_write_calc/counter/N72 ;
   wire \router/addr_calc/fft_write_calc/counter/N71 ;
   wire \router/addr_calc/fft_write_calc/counter/N70 ;
   wire \router/addr_calc/fft_write_calc/counter/N69 ;
   wire \router/addr_calc/fft_write_calc/counter/N68 ;
   wire \router/addr_calc/fft_write_calc/counter/N67 ;
   wire \router/addr_calc/fft_write_calc/counter/N66 ;
   wire \router/addr_calc/fft_write_calc/counter/N65 ;
   wire \router/addr_calc/fft_write_calc/counter/N64 ;
   wire \router/addr_calc/fft_write_calc/counter/N63 ;
   wire \router/addr_calc/fft_write_calc/counter/N62 ;
   wire \router/addr_calc/fft_write_calc/counter/N61 ;
   wire \router/addr_calc/fft_write_calc/counter/N60 ;
   wire \router/addr_calc/fft_write_calc/counter/N59 ;
   wire \router/addr_calc/fft_write_calc/counter/N58 ;
   wire \router/addr_calc/fft_write_calc/counter/N57 ;
   wire \router/addr_calc/fft_write_calc/counter/N56 ;
   wire \router/addr_calc/fft_write_calc/counter/N55 ;
   wire \router/addr_calc/fft_write_calc/counter/N54 ;
   wire \router/addr_calc/fft_write_calc/counter/N53 ;
   wire \router/addr_calc/fft_write_calc/counter/N52 ;
   wire \router/addr_calc/fft_write_calc/counter/N51 ;
   wire \router/addr_calc/fft_write_calc/counter/N50 ;
   wire \router/addr_calc/fft_write_calc/counter/N49 ;
   wire \router/addr_calc/fft_write_calc/counter/N48 ;
   wire \router/addr_calc/fft_write_calc/counter/N47 ;
   wire \router/addr_calc/fft_write_calc/counter/N40 ;
   wire \router/addr_calc/fft_write_calc/counter/hold ;
   wire \router/addr_calc/fir_read_calc/counter/N209 ;
   wire \router/addr_calc/fir_read_calc/counter/N208 ;
   wire \router/addr_calc/fir_read_calc/counter/N207 ;
   wire \router/addr_calc/fir_read_calc/counter/N206 ;
   wire \router/addr_calc/fir_read_calc/counter/N205 ;
   wire \router/addr_calc/fir_read_calc/counter/N204 ;
   wire \router/addr_calc/fir_read_calc/counter/N203 ;
   wire \router/addr_calc/fir_read_calc/counter/N202 ;
   wire \router/addr_calc/fir_read_calc/counter/N201 ;
   wire \router/addr_calc/fir_read_calc/counter/N200 ;
   wire \router/addr_calc/fir_read_calc/counter/N199 ;
   wire \router/addr_calc/fir_read_calc/counter/N198 ;
   wire \router/addr_calc/fir_read_calc/counter/N197 ;
   wire \router/addr_calc/fir_read_calc/counter/N196 ;
   wire \router/addr_calc/fir_read_calc/counter/N195 ;
   wire \router/addr_calc/fir_read_calc/counter/N194 ;
   wire \router/addr_calc/fir_read_calc/counter/N193 ;
   wire \router/addr_calc/fir_read_calc/counter/N192 ;
   wire \router/addr_calc/fir_read_calc/counter/N191 ;
   wire \router/addr_calc/fir_read_calc/counter/N190 ;
   wire \router/addr_calc/fir_read_calc/counter/N189 ;
   wire \router/addr_calc/fir_read_calc/counter/N188 ;
   wire \router/addr_calc/fir_read_calc/counter/N187 ;
   wire \router/addr_calc/fir_read_calc/counter/N186 ;
   wire \router/addr_calc/fir_read_calc/counter/N185 ;
   wire \router/addr_calc/fir_read_calc/counter/N184 ;
   wire \router/addr_calc/fir_read_calc/counter/N183 ;
   wire \router/addr_calc/fir_read_calc/counter/N182 ;
   wire \router/addr_calc/fir_read_calc/counter/N181 ;
   wire \router/addr_calc/fir_read_calc/counter/N180 ;
   wire \router/addr_calc/fir_read_calc/counter/N179 ;
   wire \router/addr_calc/fir_read_calc/counter/N178 ;
   wire \router/addr_calc/fir_read_calc/counter/N77 ;
   wire \router/addr_calc/fir_read_calc/counter/N76 ;
   wire \router/addr_calc/fir_read_calc/counter/N75 ;
   wire \router/addr_calc/fir_read_calc/counter/N74 ;
   wire \router/addr_calc/fir_read_calc/counter/N73 ;
   wire \router/addr_calc/fir_read_calc/counter/N72 ;
   wire \router/addr_calc/fir_read_calc/counter/N71 ;
   wire \router/addr_calc/fir_read_calc/counter/N70 ;
   wire \router/addr_calc/fir_read_calc/counter/N69 ;
   wire \router/addr_calc/fir_read_calc/counter/N68 ;
   wire \router/addr_calc/fir_read_calc/counter/N67 ;
   wire \router/addr_calc/fir_read_calc/counter/N66 ;
   wire \router/addr_calc/fir_read_calc/counter/N65 ;
   wire \router/addr_calc/fir_read_calc/counter/N64 ;
   wire \router/addr_calc/fir_read_calc/counter/N63 ;
   wire \router/addr_calc/fir_read_calc/counter/N62 ;
   wire \router/addr_calc/fir_read_calc/counter/N61 ;
   wire \router/addr_calc/fir_read_calc/counter/N60 ;
   wire \router/addr_calc/fir_read_calc/counter/N59 ;
   wire \router/addr_calc/fir_read_calc/counter/N58 ;
   wire \router/addr_calc/fir_read_calc/counter/N57 ;
   wire \router/addr_calc/fir_read_calc/counter/N56 ;
   wire \router/addr_calc/fir_read_calc/counter/N55 ;
   wire \router/addr_calc/fir_read_calc/counter/N54 ;
   wire \router/addr_calc/fir_read_calc/counter/N53 ;
   wire \router/addr_calc/fir_read_calc/counter/N52 ;
   wire \router/addr_calc/fir_read_calc/counter/N51 ;
   wire \router/addr_calc/fir_read_calc/counter/N50 ;
   wire \router/addr_calc/fir_read_calc/counter/N49 ;
   wire \router/addr_calc/fir_read_calc/counter/N48 ;
   wire \router/addr_calc/fir_read_calc/counter/N47 ;
   wire \router/addr_calc/fir_read_calc/counter/N40 ;
   wire \router/addr_calc/fir_read_calc/counter/hold ;
   wire \router/addr_calc/fir_write_calc/counter/N209 ;
   wire \router/addr_calc/fir_write_calc/counter/N208 ;
   wire \router/addr_calc/fir_write_calc/counter/N207 ;
   wire \router/addr_calc/fir_write_calc/counter/N206 ;
   wire \router/addr_calc/fir_write_calc/counter/N205 ;
   wire \router/addr_calc/fir_write_calc/counter/N204 ;
   wire \router/addr_calc/fir_write_calc/counter/N203 ;
   wire \router/addr_calc/fir_write_calc/counter/N202 ;
   wire \router/addr_calc/fir_write_calc/counter/N201 ;
   wire \router/addr_calc/fir_write_calc/counter/N200 ;
   wire \router/addr_calc/fir_write_calc/counter/N199 ;
   wire \router/addr_calc/fir_write_calc/counter/N198 ;
   wire \router/addr_calc/fir_write_calc/counter/N197 ;
   wire \router/addr_calc/fir_write_calc/counter/N196 ;
   wire \router/addr_calc/fir_write_calc/counter/N195 ;
   wire \router/addr_calc/fir_write_calc/counter/N194 ;
   wire \router/addr_calc/fir_write_calc/counter/N193 ;
   wire \router/addr_calc/fir_write_calc/counter/N192 ;
   wire \router/addr_calc/fir_write_calc/counter/N191 ;
   wire \router/addr_calc/fir_write_calc/counter/N190 ;
   wire \router/addr_calc/fir_write_calc/counter/N189 ;
   wire \router/addr_calc/fir_write_calc/counter/N188 ;
   wire \router/addr_calc/fir_write_calc/counter/N187 ;
   wire \router/addr_calc/fir_write_calc/counter/N186 ;
   wire \router/addr_calc/fir_write_calc/counter/N185 ;
   wire \router/addr_calc/fir_write_calc/counter/N184 ;
   wire \router/addr_calc/fir_write_calc/counter/N183 ;
   wire \router/addr_calc/fir_write_calc/counter/N182 ;
   wire \router/addr_calc/fir_write_calc/counter/N181 ;
   wire \router/addr_calc/fir_write_calc/counter/N180 ;
   wire \router/addr_calc/fir_write_calc/counter/N179 ;
   wire \router/addr_calc/fir_write_calc/counter/N178 ;
   wire \router/addr_calc/fir_write_calc/counter/N77 ;
   wire \router/addr_calc/fir_write_calc/counter/N76 ;
   wire \router/addr_calc/fir_write_calc/counter/N75 ;
   wire \router/addr_calc/fir_write_calc/counter/N74 ;
   wire \router/addr_calc/fir_write_calc/counter/N73 ;
   wire \router/addr_calc/fir_write_calc/counter/N72 ;
   wire \router/addr_calc/fir_write_calc/counter/N71 ;
   wire \router/addr_calc/fir_write_calc/counter/N70 ;
   wire \router/addr_calc/fir_write_calc/counter/N69 ;
   wire \router/addr_calc/fir_write_calc/counter/N68 ;
   wire \router/addr_calc/fir_write_calc/counter/N67 ;
   wire \router/addr_calc/fir_write_calc/counter/N66 ;
   wire \router/addr_calc/fir_write_calc/counter/N65 ;
   wire \router/addr_calc/fir_write_calc/counter/N64 ;
   wire \router/addr_calc/fir_write_calc/counter/N63 ;
   wire \router/addr_calc/fir_write_calc/counter/N62 ;
   wire \router/addr_calc/fir_write_calc/counter/N61 ;
   wire \router/addr_calc/fir_write_calc/counter/N60 ;
   wire \router/addr_calc/fir_write_calc/counter/N59 ;
   wire \router/addr_calc/fir_write_calc/counter/N58 ;
   wire \router/addr_calc/fir_write_calc/counter/N57 ;
   wire \router/addr_calc/fir_write_calc/counter/N56 ;
   wire \router/addr_calc/fir_write_calc/counter/N55 ;
   wire \router/addr_calc/fir_write_calc/counter/N54 ;
   wire \router/addr_calc/fir_write_calc/counter/N53 ;
   wire \router/addr_calc/fir_write_calc/counter/N52 ;
   wire \router/addr_calc/fir_write_calc/counter/N51 ;
   wire \router/addr_calc/fir_write_calc/counter/N50 ;
   wire \router/addr_calc/fir_write_calc/counter/N49 ;
   wire \router/addr_calc/fir_write_calc/counter/N48 ;
   wire \router/addr_calc/fir_write_calc/counter/N47 ;
   wire \router/addr_calc/fir_write_calc/counter/N40 ;
   wire \router/addr_calc/fir_write_calc/counter/hold ;
   wire \router/addr_calc/iir_read_calc/counter/N40 ;
   wire \router/addr_calc/iir_write_calc/counter/N212 ;
   wire \router/addr_calc/iir_write_calc/counter/N209 ;
   wire \router/addr_calc/iir_write_calc/counter/N208 ;
   wire \router/addr_calc/iir_write_calc/counter/N207 ;
   wire \router/addr_calc/iir_write_calc/counter/N206 ;
   wire \router/addr_calc/iir_write_calc/counter/N205 ;
   wire \router/addr_calc/iir_write_calc/counter/N204 ;
   wire \router/addr_calc/iir_write_calc/counter/N203 ;
   wire \router/addr_calc/iir_write_calc/counter/N202 ;
   wire \router/addr_calc/iir_write_calc/counter/N201 ;
   wire \router/addr_calc/iir_write_calc/counter/N200 ;
   wire \router/addr_calc/iir_write_calc/counter/N199 ;
   wire \router/addr_calc/iir_write_calc/counter/N198 ;
   wire \router/addr_calc/iir_write_calc/counter/N197 ;
   wire \router/addr_calc/iir_write_calc/counter/N196 ;
   wire \router/addr_calc/iir_write_calc/counter/N195 ;
   wire \router/addr_calc/iir_write_calc/counter/N194 ;
   wire \router/addr_calc/iir_write_calc/counter/N193 ;
   wire \router/addr_calc/iir_write_calc/counter/N192 ;
   wire \router/addr_calc/iir_write_calc/counter/N191 ;
   wire \router/addr_calc/iir_write_calc/counter/N190 ;
   wire \router/addr_calc/iir_write_calc/counter/N189 ;
   wire \router/addr_calc/iir_write_calc/counter/N188 ;
   wire \router/addr_calc/iir_write_calc/counter/N187 ;
   wire \router/addr_calc/iir_write_calc/counter/N186 ;
   wire \router/addr_calc/iir_write_calc/counter/N185 ;
   wire \router/addr_calc/iir_write_calc/counter/N184 ;
   wire \router/addr_calc/iir_write_calc/counter/N183 ;
   wire \router/addr_calc/iir_write_calc/counter/N182 ;
   wire \router/addr_calc/iir_write_calc/counter/N181 ;
   wire \router/addr_calc/iir_write_calc/counter/N180 ;
   wire \router/addr_calc/iir_write_calc/counter/N179 ;
   wire \router/addr_calc/iir_write_calc/counter/N178 ;
   wire \router/addr_calc/iir_write_calc/counter/N76 ;
   wire \router/addr_calc/iir_write_calc/counter/N75 ;
   wire \router/addr_calc/iir_write_calc/counter/N74 ;
   wire \router/addr_calc/iir_write_calc/counter/N73 ;
   wire \router/addr_calc/iir_write_calc/counter/N72 ;
   wire \router/addr_calc/iir_write_calc/counter/N71 ;
   wire \router/addr_calc/iir_write_calc/counter/N70 ;
   wire \router/addr_calc/iir_write_calc/counter/N69 ;
   wire \router/addr_calc/iir_write_calc/counter/N68 ;
   wire \router/addr_calc/iir_write_calc/counter/N67 ;
   wire \router/addr_calc/iir_write_calc/counter/N66 ;
   wire \router/addr_calc/iir_write_calc/counter/N65 ;
   wire \router/addr_calc/iir_write_calc/counter/N64 ;
   wire \router/addr_calc/iir_write_calc/counter/N63 ;
   wire \router/addr_calc/iir_write_calc/counter/N62 ;
   wire \router/addr_calc/iir_write_calc/counter/N61 ;
   wire \router/addr_calc/iir_write_calc/counter/N60 ;
   wire \router/addr_calc/iir_write_calc/counter/N59 ;
   wire \router/addr_calc/iir_write_calc/counter/N58 ;
   wire \router/addr_calc/iir_write_calc/counter/N57 ;
   wire \router/addr_calc/iir_write_calc/counter/N56 ;
   wire \router/addr_calc/iir_write_calc/counter/N55 ;
   wire \router/addr_calc/iir_write_calc/counter/N54 ;
   wire \router/addr_calc/iir_write_calc/counter/N53 ;
   wire \router/addr_calc/iir_write_calc/counter/N52 ;
   wire \router/addr_calc/iir_write_calc/counter/N51 ;
   wire \router/addr_calc/iir_write_calc/counter/N50 ;
   wire \router/addr_calc/iir_write_calc/counter/N49 ;
   wire \router/addr_calc/iir_write_calc/counter/N48 ;
   wire \router/addr_calc/iir_write_calc/counter/N47 ;
   wire \router/addr_calc/iir_write_calc/counter/N40 ;
   wire \router/addr_calc/iir_write_calc/counter/hold ;
   wire \fifo_to_fir/fifo_cell0/reg_ptok/N29 ;
   wire \fifo_to_fft/fifo_cell0/reg_ptok/N29 ;
   wire \fifo_from_fir/fifo_cell0/reg_ptok/N29 ;
   wire \fifo_from_fft/fifo_cell0/reg_ptok/N29 ;
   wire \fifo_from_fir/fifo_cell0/data_out/N9 ;
   wire \fifo_from_fft/fifo_cell0/data_out/N9 ;
   wire n137;
   wire n521;
   wire n585;
   wire n649;
   wire n713;
   wire n777;
   wire n841;
   wire n905;
   wire n969;
   wire n1033;
   wire n1097;
   wire n1161;
   wire n1225;
   wire n1289;
   wire n1353;
   wire n1417;
   wire n1481;
   wire n1545;
   wire n1609;
   wire n1673;
   wire n1737;
   wire n1801;
   wire n1865;
   wire n1929;
   wire n1993;
   wire n2057;
   wire n2121;
   wire n2185;
   wire n2249;
   wire n2313;
   wire n2377;
   wire n2441;
   wire n2505;
   wire n2569;
   wire n2633;
   wire n2634;
   wire n2804;
   wire n2807;
   wire n2810;
   wire n2813;
   wire n2816;
   wire n2819;
   wire n2822;
   wire n2825;
   wire n2828;
   wire n2831;
   wire n2834;
   wire n2837;
   wire n2840;
   wire n2843;
   wire n2848;
   wire n2852;
   wire n2855;
   wire n2858;
   wire n2861;
   wire n2864;
   wire n2867;
   wire n2870;
   wire n2873;
   wire n2876;
   wire n2879;
   wire n2882;
   wire n2885;
   wire n2888;
   wire n2891;
   wire n3440;
   wire n3455;
   wire n3456;
   wire n3458;
   wire n3463;
   wire n3465;
   wire n3467;
   wire n3468;
   wire n3469;
   wire n3470;
   wire n3471;
   wire n3472;
   wire n3473;
   wire n3474;
   wire n3476;
   wire n3477;
   wire n3478;
   wire n3479;
   wire n3480;
   wire n3481;
   wire n3482;
   wire n3483;
   wire n3484;
   wire n3486;
   wire n3487;
   wire n3488;
   wire n3489;
   wire n3490;
   wire n3491;
   wire n3492;
   wire n3493;
   wire n3494;
   wire n3495;
   wire n3496;
   wire n3497;
   wire n3498;
   wire n3499;
   wire n3500;
   wire n3501;
   wire n3502;
   wire n3503;
   wire n3504;
   wire n3505;
   wire n3506;
   wire n3507;
   wire n3508;
   wire n3509;
   wire n3510;
   wire n3511;
   wire n3512;
   wire n3513;
   wire n3514;
   wire n3515;
   wire n3516;
   wire n3517;
   wire n3518;
   wire n3519;
   wire n3520;
   wire n3521;
   wire n3522;
   wire n3523;
   wire n3524;
   wire n3525;
   wire n3526;
   wire n3527;
   wire n3528;
   wire n3529;
   wire n3530;
   wire n3531;
   wire n3532;
   wire n3533;
   wire n3534;
   wire n3535;
   wire n3536;
   wire n3537;
   wire n3538;
   wire n3539;
   wire n3540;
   wire n3541;
   wire n3542;
   wire n3543;
   wire n3544;
   wire n3545;
   wire n3546;
   wire n3547;
   wire n3548;
   wire n3549;
   wire n3550;
   wire n3551;
   wire n3552;
   wire n3553;
   wire n3554;
   wire n3555;
   wire n3556;
   wire n3557;
   wire n3558;
   wire n3559;
   wire n3560;
   wire n3561;
   wire n3562;
   wire n3563;
   wire n3564;
   wire n3565;
   wire n3566;
   wire n3567;
   wire n3568;
   wire n3569;
   wire n3570;
   wire n3571;
   wire n3572;
   wire n3573;
   wire n3574;
   wire n3575;
   wire n3576;
   wire n3577;
   wire n3578;
   wire n3579;
   wire n3580;
   wire n3581;
   wire n3582;
   wire n3583;
   wire n3584;
   wire n3585;
   wire n3586;
   wire n3587;
   wire n3588;
   wire n3589;
   wire n3590;
   wire n3591;
   wire n3592;
   wire n3593;
   wire n3594;
   wire n3595;
   wire n3596;
   wire n3597;
   wire n3598;
   wire n3599;
   wire n3600;
   wire n3601;
   wire n3602;
   wire n3603;
   wire n3604;
   wire n3605;
   wire n3606;
   wire n3607;
   wire n3608;
   wire n3609;
   wire n3610;
   wire n3611;
   wire n3612;
   wire n3613;
   wire n3614;
   wire n3615;
   wire n3616;
   wire n3617;
   wire n3618;
   wire n3619;
   wire n3620;
   wire n3621;
   wire n3622;
   wire n3623;
   wire n3624;
   wire n3625;
   wire n3626;
   wire n3627;
   wire n3628;
   wire n3629;
   wire n3630;
   wire n3631;
   wire n3632;
   wire n3633;
   wire n3634;
   wire n3635;
   wire n3636;
   wire n3637;
   wire n3638;
   wire n3639;
   wire n3640;
   wire n3641;
   wire n3642;
   wire n3643;
   wire n3644;
   wire n3645;
   wire n3646;
   wire n3647;
   wire n3648;
   wire n3649;
   wire n3650;
   wire n3651;
   wire n3652;
   wire n3653;
   wire n3654;
   wire n3655;
   wire n3656;
   wire n3657;
   wire n3658;
   wire n3659;
   wire n3660;
   wire n3661;
   wire n3662;
   wire n3663;
   wire n3664;
   wire n3665;
   wire n3666;
   wire n3667;
   wire n3668;
   wire n3669;
   wire n3670;
   wire n3671;
   wire n3672;
   wire n3673;
   wire n3674;
   wire n3675;
   wire n3676;
   wire n3677;
   wire n3678;
   wire n3679;
   wire n3680;
   wire n3681;
   wire n3682;
   wire n3683;
   wire n3684;
   wire n3685;
   wire n3686;
   wire n3687;
   wire n3688;
   wire n3689;
   wire n3690;
   wire n3691;
   wire n3692;
   wire n3693;
   wire n3694;
   wire n3695;
   wire n3696;
   wire n3697;
   wire n3698;
   wire n3699;
   wire n3700;
   wire n3701;
   wire n3702;
   wire n3703;
   wire n3704;
   wire n3705;
   wire n3706;
   wire n3707;
   wire n3708;
   wire n3709;
   wire n3710;
   wire n3712;
   wire n3713;
   wire n3714;
   wire n3715;
   wire n3716;
   wire n3717;
   wire n3719;
   wire n3720;
   wire n3721;
   wire n3722;
   wire n3723;
   wire n3724;
   wire n3725;
   wire n3726;
   wire n3727;
   wire n3728;
   wire n3729;
   wire n3730;
   wire n3731;
   wire n3732;
   wire n3733;
   wire n3734;
   wire n3735;
   wire n3736;
   wire n3737;
   wire n3738;
   wire n3739;
   wire n3740;
   wire n3741;
   wire n3742;
   wire n3743;
   wire n3744;
   wire n3745;
   wire n3746;
   wire n3747;
   wire n3748;
   wire n3749;
   wire n3750;
   wire n3751;
   wire n3752;
   wire n3753;
   wire n3754;
   wire n3755;
   wire n3756;
   wire n3757;
   wire n3758;
   wire n3760;
   wire n3763;
   wire n3764;
   wire n3767;
   wire n3768;
   wire n3769;
   wire n3771;
   wire n3772;
   wire n3774;
   wire n3776;
   wire n3777;
   wire n3778;
   wire n3780;
   wire n3783;
   wire n3784;
   wire n3787;
   wire n3788;
   wire n3789;
   wire n3791;
   wire n3792;
   wire n3794;
   wire n3796;
   wire n3797;
   wire n3798;
   wire n3800;
   wire n3803;
   wire n3804;
   wire n3807;
   wire n3808;
   wire n3809;
   wire n3811;
   wire n3814;
   wire n3815;
   wire n3818;
   wire n3819;
   wire n3820;
   wire n3823;
   wire n3824;
   wire n3825;
   wire n3826;
   wire n3827;
   wire n3828;
   wire n3829;
   wire n3830;
   wire n3831;
   wire n3832;
   wire n3833;
   wire n3834;
   wire n3835;
   wire n3837;
   wire n3838;
   wire n3839;
   wire n3840;
   wire n3841;
   wire n3842;
   wire n3843;
   wire n3844;
   wire n3845;
   wire n3846;
   wire n3847;
   wire n3848;
   wire n3849;
   wire n3850;
   wire n3851;
   wire n3854;
   wire n3855;
   wire n3856;
   wire n3857;
   wire n3858;
   wire n3859;
   wire n3860;
   wire n3861;
   wire n3862;
   wire n3863;
   wire n3864;
   wire n3865;
   wire n3866;
   wire n3867;
   wire n3868;
   wire n3869;
   wire n3870;
   wire n3871;
   wire n3872;
   wire n3873;
   wire n3874;
   wire n3875;
   wire n3876;
   wire n3877;
   wire n3878;
   wire n3879;
   wire n3880;
   wire n3881;
   wire n3883;
   wire n3884;
   wire n3885;
   wire n3886;
   wire n3887;
   wire n3888;
   wire n3889;
   wire n3890;
   wire n3891;
   wire n3892;
   wire n3893;
   wire n3894;
   wire n3895;
   wire n3896;
   wire n3897;
   wire n3898;
   wire n3899;
   wire n3900;
   wire n3901;
   wire n3902;
   wire n3903;
   wire n3904;
   wire n3905;
   wire n3906;
   wire n3907;
   wire n3908;
   wire n3909;
   wire n3910;
   wire n3911;
   wire n3912;
   wire n3913;
   wire n3914;
   wire n3915;
   wire n3916;
   wire n3917;
   wire n3918;
   wire n3919;
   wire n3920;
   wire n3921;
   wire n3922;
   wire n3923;
   wire n3924;
   wire n3925;
   wire n3926;
   wire n3927;
   wire n3928;
   wire n3929;
   wire n3930;
   wire n3931;
   wire n3932;
   wire n3933;
   wire n3934;
   wire n3935;
   wire n3936;
   wire n3937;
   wire n3938;
   wire n3939;
   wire n3940;
   wire n3941;
   wire n3942;
   wire n3943;
   wire n3944;
   wire n3945;
   wire n3946;
   wire n3947;
   wire n3948;
   wire n3949;
   wire n3950;
   wire n3951;
   wire n3952;
   wire n3953;
   wire n3954;
   wire n3955;
   wire n3956;
   wire n3957;
   wire n3958;
   wire n3959;
   wire n3960;
   wire n3961;
   wire n3962;
   wire n3963;
   wire n3964;
   wire n3965;
   wire n3966;
   wire n3967;
   wire n3968;
   wire n3969;
   wire n3970;
   wire n3971;
   wire n3972;
   wire n3973;
   wire n3974;
   wire n3975;
   wire n3976;
   wire n3977;
   wire n3978;
   wire n3979;
   wire n3980;
   wire n3981;
   wire n3982;
   wire n3983;
   wire n3984;
   wire n3985;
   wire n3986;
   wire n3987;
   wire n3988;
   wire n3989;
   wire n3990;
   wire n3991;
   wire n3992;
   wire n3993;
   wire n3994;
   wire n3995;
   wire n3996;
   wire n3997;
   wire n3998;
   wire n3999;
   wire n4000;
   wire n4001;
   wire n4003;
   wire n4004;
   wire n4005;
   wire n4006;
   wire n4009;
   wire n4023;
   wire n4025;
   wire n4026;
   wire n4029;
   wire n4030;
   wire n4031;
   wire n4032;
   wire n4033;
   wire n4034;
   wire n4035;
   wire n4036;
   wire n4037;
   wire n4038;
   wire n4039;
   wire n4040;
   wire n4041;
   wire n4042;
   wire n4043;
   wire n4044;
   wire n4045;
   wire n4046;
   wire n4047;
   wire n4048;
   wire n4049;
   wire n4050;
   wire n4051;
   wire n4052;
   wire n4053;
   wire n4054;
   wire n4055;
   wire n4056;
   wire n4057;
   wire n4058;
   wire n4059;
   wire n4060;
   wire n4061;
   wire n4062;
   wire n4063;
   wire n4064;
   wire n4065;
   wire n4066;
   wire n4067;
   wire n4068;
   wire n4069;
   wire n4070;
   wire n4071;
   wire n4072;
   wire n4073;
   wire n4074;
   wire n4075;
   wire n4076;
   wire n4077;
   wire n4078;
   wire n4079;
   wire n4080;
   wire n4081;
   wire n4082;
   wire n4083;
   wire n4084;
   wire n4085;
   wire n4086;
   wire n4087;
   wire n4088;
   wire n4089;
   wire n4090;
   wire n4091;
   wire n4092;
   wire n4093;
   wire n4094;
   wire n4095;
   wire n4096;
   wire n4097;
   wire n4098;
   wire n4099;
   wire n4100;
   wire n4101;
   wire n4102;
   wire n4103;
   wire n4104;
   wire n4105;
   wire n4106;
   wire n4107;
   wire n4108;
   wire n4109;
   wire n4110;
   wire n4111;
   wire n4112;
   wire n4113;
   wire n4114;
   wire n4115;
   wire n4116;
   wire n4117;
   wire n4118;
   wire n4119;
   wire n4120;
   wire n4121;
   wire n4122;
   wire n4123;
   wire n4124;
   wire n4125;
   wire n4126;
   wire n4127;
   wire n4128;
   wire n4129;
   wire n4130;
   wire n4131;
   wire n4132;
   wire n4133;
   wire n4134;
   wire n4135;
   wire n4136;
   wire n4137;
   wire n4138;
   wire n4139;
   wire n4140;
   wire n4141;
   wire n4142;
   wire n4143;
   wire n4144;
   wire n4145;
   wire n4146;
   wire n4147;
   wire n4148;
   wire n4149;
   wire n4150;
   wire n4151;
   wire n4152;
   wire n4153;
   wire n4154;
   wire n4155;
   wire n4156;
   wire n4157;
   wire n4158;
   wire n4159;
   wire n4160;
   wire n4161;
   wire n4162;
   wire n4163;
   wire n4164;
   wire n4165;
   wire n4166;
   wire n4167;
   wire n4168;
   wire n4169;
   wire n4170;
   wire n4171;
   wire n4172;
   wire n4173;
   wire n4174;
   wire n4175;
   wire n4176;
   wire n4178;
   wire n4179;
   wire n4180;
   wire n4181;
   wire n4184;
   wire n4198;
   wire n4200;
   wire n4201;
   wire n4202;
   wire n4203;
   wire n4204;
   wire n4205;
   wire n4207;
   wire n4311;
   wire n4441;
   wire n4442;
   wire n4443;
   wire n4444;
   wire n4445;
   wire n4449;
   wire n4450;
   wire n4451;
   wire n4452;
   wire n4453;
   wire n4454;
   wire n4455;
   wire n4456;
   wire n4457;
   wire n4458;
   wire n4459;
   wire n4460;
   wire n4461;
   wire n4462;
   wire n4463;
   wire n4464;
   wire n4465;
   wire n4466;
   wire n4467;
   wire n4468;
   wire n4469;
   wire n4470;
   wire n4471;
   wire n4472;
   wire n4473;
   wire n4474;
   wire n4475;
   wire n4476;
   wire n4477;
   wire n4478;
   wire n4479;
   wire n4480;
   wire n4481;
   wire n4482;
   wire n4483;
   wire n4484;
   wire n4485;
   wire n4486;
   wire n4487;
   wire n4488;
   wire n4489;
   wire n4490;
   wire n4491;
   wire n4492;
   wire n4493;
   wire n4494;
   wire n4495;
   wire n4496;
   wire n4497;
   wire n4498;
   wire n4499;
   wire n4500;
   wire n4502;
   wire n4503;
   wire n4504;
   wire n4505;
   wire n4506;
   wire n4507;
   wire n4508;
   wire n4509;
   wire n4510;
   wire n4511;
   wire n4512;
   wire n4513;
   wire n4514;
   wire n4515;
   wire n4516;
   wire n4517;
   wire n4518;
   wire n4519;
   wire n4520;
   wire n4521;
   wire n4522;
   wire n4523;
   wire n4524;
   wire n4525;
   wire n4526;
   wire n4527;
   wire n4528;
   wire n4529;
   wire n4530;
   wire n4531;
   wire n4532;
   wire n4533;
   wire n4534;
   wire n4535;
   wire n4536;
   wire n4537;
   wire n4538;
   wire n4539;
   wire n4540;
   wire n4541;
   wire n4542;
   wire n4543;
   wire n4544;
   wire n4545;
   wire n4546;
   wire n4547;
   wire n4548;
   wire n4549;
   wire n4550;
   wire n4551;
   wire n4552;
   wire n4553;
   wire n4554;
   wire n4555;
   wire n4556;
   wire n4557;
   wire n4558;
   wire n4559;
   wire n4560;
   wire n4561;
   wire n4562;
   wire n4563;
   wire n4564;
   wire n4565;
   wire n4566;
   wire n4568;
   wire n4569;
   wire n4570;
   wire n4571;
   wire n4572;
   wire n4573;
   wire n4574;
   wire n4575;
   wire n4576;
   wire n4577;
   wire n4578;
   wire n4579;
   wire n4580;
   wire n4595;
   wire n4597;
   wire n4598;
   wire n4599;
   wire n4600;
   wire n4601;
   wire n4602;
   wire n4603;
   wire n4604;
   wire n4605;
   wire n4606;
   wire n4607;
   wire n4608;
   wire n4609;
   wire n4610;
   wire n4611;
   wire n4612;
   wire n4613;
   wire n4614;
   wire n4615;
   wire n4616;
   wire n4617;
   wire n4618;
   wire n4619;
   wire n4620;
   wire n4621;
   wire n4622;
   wire n4623;
   wire n4624;
   wire n4625;
   wire n4626;
   wire n4627;
   wire n4628;
   wire n4629;
   wire n4630;
   wire n4631;
   wire n4632;
   wire n4633;
   wire n4634;
   wire n4635;
   wire n4636;
   wire n4637;
   wire n4638;
   wire n4639;
   wire n4640;
   wire n4641;
   wire n4643;
   wire n4644;
   wire n4645;
   wire n4646;
   wire n4647;
   wire n4648;
   wire n4649;
   wire n4650;
   wire n4651;
   wire n4652;
   wire n4653;
   wire n4654;
   wire n4655;
   wire n4656;
   wire n4657;
   wire n4658;
   wire n4659;
   wire n4660;
   wire n4661;
   wire n4662;
   wire n4663;
   wire n4664;
   wire n4665;
   wire n4666;
   wire n4667;
   wire n4668;
   wire n4669;
   wire n4670;
   wire n4671;
   wire n4672;
   wire n4673;
   wire n4674;
   wire n4675;
   wire n4676;
   wire n4677;
   wire n4678;
   wire n4679;
   wire n4680;
   wire n4681;
   wire n4682;
   wire n4683;
   wire n4684;
   wire n4685;
   wire n4686;
   wire n4688;
   wire n4689;
   wire n4690;
   wire n4691;
   wire n4692;
   wire n4693;
   wire n4694;
   wire n4695;
   wire n4696;
   wire n4697;
   wire n4698;
   wire n4699;
   wire n4700;
   wire n4701;
   wire n4702;
   wire n4703;
   wire n4704;
   wire n4705;
   wire n4706;
   wire n4707;
   wire n4708;
   wire n4709;
   wire n4710;
   wire n4711;
   wire n4712;
   wire n4713;
   wire n4714;
   wire n4715;
   wire n4716;
   wire n4717;
   wire n4718;
   wire n4719;
   wire n4720;
   wire n4721;
   wire n4722;
   wire n4723;
   wire n4724;
   wire n4725;
   wire n4726;
   wire n4727;
   wire n4728;
   wire n4729;
   wire n4730;
   wire n4731;
   wire n4732;
   wire n4733;
   wire n4734;
   wire n4735;
   wire n4736;
   wire n4737;
   wire n4738;
   wire n4739;
   wire n4740;
   wire n4741;
   wire n4742;
   wire n4743;
   wire n4744;
   wire n4745;
   wire n4746;
   wire n4747;
   wire n4748;
   wire n4749;
   wire n4750;
   wire n4751;
   wire n4752;
   wire n4754;
   wire n4755;
   wire n4756;
   wire n4757;
   wire n4758;
   wire n4759;
   wire n4760;
   wire n4761;
   wire n4762;
   wire n4763;
   wire n4764;
   wire n4765;
   wire n4766;
   wire n4781;
   wire n4783;
   wire n4784;
   wire n4785;
   wire n4786;
   wire n4787;
   wire n4788;
   wire n4789;
   wire n4790;
   wire n4791;
   wire n4792;
   wire n4793;
   wire n4794;
   wire n4795;
   wire n4796;
   wire n4797;
   wire n4798;
   wire n4799;
   wire n4800;
   wire n4801;
   wire n4802;
   wire n4803;
   wire n4804;
   wire n4805;
   wire n4806;
   wire n4807;
   wire n4808;
   wire n4809;
   wire n4810;
   wire n4811;
   wire n4812;
   wire n4813;
   wire n4814;
   wire n4815;
   wire n4816;
   wire n4817;
   wire n4818;
   wire n4819;
   wire n4820;
   wire n4821;
   wire n4822;
   wire n4823;
   wire n4824;
   wire n4825;
   wire n4826;
   wire n4827;
   wire n4829;
   wire n4830;
   wire n4832;
   wire n4840;
   wire n4841;
   wire n5191;
   wire n5193;
   wire n5196;
   wire n5197;
   wire n5198;
   wire n5199;
   wire n5202;
   wire n5203;
   wire n5206;
   wire n5207;
   wire n5208;
   wire n5213;
   wire n5214;
   wire n5215;
   wire n5216;
   wire n5217;
   wire n5218;
   wire n5219;
   wire n5220;
   wire n5221;
   wire n5222;
   wire n5223;
   wire n5224;
   wire n5225;
   wire n5226;
   wire n5233;
   wire n5240;
   wire n5243;
   wire n5244;
   wire n5246;
   wire n5248;
   wire n5249;
   wire n5250;
   wire n5255;
   wire n5256;
   wire n5257;
   wire n5258;
   wire n5259;
   wire n5260;
   wire n5261;
   wire n5262;
   wire n5263;
   wire n5264;
   wire n5265;
   wire n5266;
   wire n5267;
   wire n5268;
   wire n5274;
   wire n5275;
   wire n5276;
   wire n5277;
   wire n5278;
   wire n5279;
   wire n5281;
   wire n5282;
   wire n5283;
   wire n5284;
   wire n5285;
   wire n5286;
   wire n5287;
   wire n5288;
   wire n5312;
   wire n5313;
   wire n5314;
   wire n5315;
   wire n5316;
   wire n5317;
   wire n5318;
   wire n5320;
   wire n5321;
   wire n5322;
   wire n5323;
   wire n5324;
   wire n5326;
   wire n5327;
   wire n5346;
   wire n5351;
   wire n5352;
   wire n5353;
   wire n5354;
   wire n5355;
   wire n5356;
   wire n5357;
   wire n5358;
   wire n5359;
   wire n5360;
   wire n5361;
   wire n5362;
   wire n5363;
   wire n5364;
   wire n5365;
   wire n5366;
   wire n5367;
   wire n5368;
   wire n5369;
   wire n5370;
   wire n5371;
   wire n5372;
   wire n5373;
   wire n5374;
   wire n5375;
   wire n5376;
   wire n5377;
   wire n5378;
   wire n5379;
   wire n5380;
   wire n5381;
   wire n5382;
   wire n5383;
   wire n5384;
   wire n5385;
   wire n5386;
   wire n5387;
   wire n5388;
   wire n5389;
   wire n5390;
   wire n5391;
   wire n5392;
   wire n5393;
   wire n5394;
   wire n5395;
   wire n5396;
   wire n5397;
   wire n5398;
   wire n5399;
   wire n5400;
   wire n5401;
   wire n5402;
   wire n5403;
   wire n5404;
   wire n5405;
   wire n5406;
   wire n5407;
   wire n5408;
   wire n5409;
   wire n5410;
   wire n5411;
   wire n5412;
   wire n5413;
   wire n5414;
   wire n5415;
   wire n5416;
   wire n5417;
   wire n5418;
   wire n5419;
   wire n5420;
   wire n5421;
   wire n5422;
   wire n5423;
   wire n5424;
   wire n5425;
   wire n5426;
   wire n5427;
   wire n5428;
   wire n5429;
   wire n5430;
   wire n5431;
   wire n5432;
   wire n5433;
   wire n5434;
   wire n5435;
   wire n5436;
   wire n5437;
   wire n5438;
   wire n5439;
   wire n5440;
   wire n5441;
   wire n5442;
   wire n5443;
   wire n5444;
   wire n5445;
   wire n5446;
   wire n5447;
   wire n5448;
   wire n5449;
   wire n5450;
   wire n5451;
   wire n5452;
   wire n5453;
   wire n5454;
   wire n5455;
   wire n5456;
   wire n5457;
   wire n5459;
   wire n5460;
   wire n5461;
   wire n5462;
   wire n5463;
   wire n5464;
   wire n5465;
   wire n5466;
   wire n5467;
   wire n5468;
   wire n5469;
   wire n5470;
   wire n5471;
   wire n5472;
   wire n5473;
   wire n5474;
   wire n5475;
   wire n5476;
   wire n5477;
   wire n5478;
   wire n5479;
   wire n5480;
   wire n5481;
   wire n5482;
   wire n5483;
   wire n5484;
   wire n5485;
   wire n5486;
   wire n5487;
   wire n5488;
   wire n5489;
   wire n5490;
   wire n5491;
   wire n5492;
   wire n5493;
   wire n5494;
   wire n5495;
   wire n5496;
   wire n5497;
   wire n5498;
   wire n5499;
   wire n5500;
   wire n5501;
   wire n5502;
   wire n5503;
   wire n5504;
   wire n5505;
   wire n5506;
   wire n5507;
   wire n5508;
   wire n5509;
   wire n5510;
   wire n5511;
   wire n5512;
   wire n5513;
   wire n5514;
   wire n5515;
   wire n5516;
   wire n5517;
   wire n5518;
   wire n5519;
   wire n5520;
   wire n5521;
   wire n5522;
   wire n5523;
   wire n5524;
   wire n5525;
   wire n5526;
   wire n5527;
   wire n5528;
   wire n5529;
   wire n5530;
   wire n5531;
   wire n5532;
   wire n5533;
   wire n5534;
   wire n5535;
   wire n5536;
   wire n5537;
   wire n5538;
   wire n5539;
   wire n5540;
   wire n5541;
   wire n5542;
   wire n5543;
   wire n5544;
   wire n5545;
   wire n5546;
   wire n5547;
   wire n5548;
   wire n5549;
   wire n5550;
   wire n5551;
   wire n5552;
   wire n5553;
   wire n5554;
   wire n5555;
   wire n5556;
   wire n5557;
   wire n5558;
   wire n5559;
   wire n5560;
   wire n5561;
   wire n5562;
   wire n5563;
   wire n5564;
   wire n5565;
   wire n5566;
   wire n5567;
   wire n5568;
   wire n5569;
   wire n5570;
   wire n5571;
   wire n5572;
   wire n5573;
   wire n5574;
   wire n5575;
   wire n5576;
   wire n5577;
   wire n5578;
   wire n5579;
   wire n5580;
   wire n5581;
   wire n5582;
   wire n5583;
   wire n5584;
   wire n5585;
   wire n5586;
   wire n5587;
   wire n5588;
   wire n5589;
   wire n5590;
   wire n5591;
   wire n5592;
   wire n5593;
   wire n5594;
   wire n5595;
   wire n5596;
   wire n5597;
   wire n5598;
   wire n5599;
   wire n5600;
   wire n5601;
   wire n5602;
   wire n5603;
   wire n5604;
   wire n5605;
   wire n5700;
   wire n5701;
   wire n5702;
   wire n5703;
   wire n5704;
   wire n5705;
   wire n5706;
   wire n5707;
   wire n5708;
   wire n5709;
   wire n5710;
   wire n5711;
   wire n5712;
   wire n5713;
   wire n5714;
   wire n5715;
   wire n5716;
   wire n5717;
   wire n5718;
   wire n5719;
   wire n5720;
   wire n5721;
   wire n5722;
   wire n5723;
   wire n5724;
   wire n5725;
   wire n5726;
   wire n5727;
   wire n5728;
   wire n5729;
   wire n5730;
   wire n5731;
   wire n5732;
   wire n5733;
   wire n5734;
   wire n5735;
   wire n5736;
   wire n5737;
   wire n5738;
   wire n5739;
   wire n5740;
   wire n5741;
   wire n5742;
   wire n5743;
   wire n5744;
   wire n5745;
   wire n5746;
   wire n5747;
   wire n5748;
   wire n5749;
   wire n5750;
   wire n5751;
   wire n5752;
   wire n5753;
   wire n5754;
   wire n5755;
   wire n5756;
   wire n5757;
   wire n5758;
   wire n5759;
   wire n5760;
   wire n5761;
   wire n5762;
   wire n5763;
   wire n5764;
   wire n5765;
   wire n5766;
   wire n5767;
   wire n5768;
   wire n5769;
   wire n5770;
   wire n5771;
   wire n5772;
   wire n5773;
   wire n5774;
   wire n5775;
   wire n5776;
   wire n5777;
   wire n5778;
   wire n5779;
   wire n5780;
   wire n5781;
   wire n5782;
   wire n5783;
   wire n5784;
   wire n5785;
   wire n5786;
   wire n5787;
   wire n5788;
   wire n5789;
   wire n5790;
   wire n5791;
   wire n5792;
   wire n5793;
   wire n5794;
   wire n5795;
   wire n5796;
   wire n5797;
   wire n5798;
   wire n5799;
   wire n5800;
   wire n5801;
   wire n5802;
   wire n5803;
   wire n5804;
   wire n5805;
   wire n5806;
   wire n5807;
   wire n5808;
   wire n5809;
   wire n5810;
   wire n5811;
   wire n5812;
   wire n5813;
   wire n5814;
   wire n5815;
   wire n5816;
   wire n5817;
   wire n5818;
   wire n5819;
   wire n5820;
   wire n5821;
   wire n5822;
   wire n5823;
   wire n5824;
   wire n5825;
   wire n5826;
   wire n5827;
   wire n5828;
   wire n5829;
   wire n5830;
   wire n5831;
   wire n5832;
   wire n5833;
   wire n5834;
   wire n5835;
   wire n5836;
   wire n5837;
   wire n5838;
   wire n5839;
   wire n5840;
   wire n5841;
   wire n5842;
   wire n5843;
   wire n5844;
   wire n5845;
   wire n5846;
   wire n5847;
   wire n5848;
   wire n5849;
   wire n5850;
   wire n5851;
   wire n5852;
   wire n5853;
   wire n5854;
   wire n5855;
   wire n5856;
   wire n5857;
   wire n5858;
   wire n5859;
   wire n5860;
   wire n5861;
   wire n5862;
   wire n5863;
   wire n5864;
   wire n5865;
   wire n5866;
   wire n5867;
   wire n5868;
   wire n5869;
   wire n5870;
   wire n5871;
   wire n5872;
   wire n5873;
   wire n5874;
   wire n5875;
   wire n5876;
   wire n5877;
   wire n5878;
   wire n5879;
   wire n5880;
   wire n5881;
   wire n5882;
   wire n5883;
   wire n5884;
   wire n5885;
   wire n5886;
   wire n5887;
   wire n5888;
   wire n5889;
   wire n5890;
   wire n5891;
   wire n5892;
   wire n5893;
   wire n5894;
   wire n5895;
   wire n5896;
   wire n5897;
   wire n5898;
   wire n5899;
   wire n5900;
   wire n5901;
   wire n5902;
   wire n5903;
   wire n5904;
   wire n5905;
   wire n5906;
   wire n5907;
   wire n5908;
   wire n5909;
   wire n5910;
   wire n5911;
   wire n5912;
   wire n5913;
   wire n5914;
   wire n5915;
   wire n5916;
   wire n5917;
   wire n5918;
   wire n5919;
   wire n5920;
   wire n5921;
   wire n5922;
   wire n5923;
   wire n5924;
   wire n5925;
   wire n5926;
   wire n5927;
   wire n5928;
   wire n5929;
   wire n5930;
   wire n5931;
   wire n5932;
   wire n5933;
   wire n5934;
   wire n5935;
   wire n5936;
   wire n5937;
   wire n5938;
   wire n5939;
   wire n5940;
   wire n5941;
   wire n5942;
   wire n5943;
   wire n5944;
   wire n5945;
   wire n5946;
   wire n5947;
   wire n5948;
   wire n5949;
   wire n5950;
   wire n5951;
   wire n5952;
   wire n5953;
   wire n5954;
   wire n5955;
   wire n5956;
   wire n5957;
   wire n5958;
   wire n5959;
   wire n5960;
   wire n5961;
   wire n5962;
   wire n5963;
   wire n5964;
   wire n5965;
   wire n5966;
   wire n5967;
   wire n5968;
   wire n5969;
   wire n5970;
   wire n5971;
   wire n5972;
   wire n5973;
   wire n5974;
   wire n5975;
   wire n5976;
   wire n5977;
   wire n5978;
   wire n5979;
   wire n5980;
   wire n5981;
   wire n5982;
   wire n5983;
   wire n5984;
   wire n5985;
   wire n5986;
   wire n5987;
   wire n5988;
   wire n5989;
   wire n5990;
   wire n5991;
   wire n5992;
   wire n5993;
   wire n5994;
   wire n5995;
   wire n5996;
   wire n5997;
   wire n5998;
   wire n5999;
   wire n6000;
   wire n6001;
   wire n6002;
   wire n6003;
   wire n6004;
   wire n6005;
   wire n6006;
   wire n6007;
   wire n6008;
   wire n6009;
   wire n6010;
   wire n6011;
   wire n6012;
   wire n6013;
   wire n6014;
   wire n6015;
   wire n6016;
   wire n6017;
   wire n6018;
   wire n6019;
   wire n6020;
   wire n6021;
   wire n6022;
   wire n6023;
   wire n6024;
   wire n6025;
   wire n6026;
   wire n6027;
   wire n6028;
   wire n6029;
   wire n6030;
   wire n6031;
   wire n6032;
   wire n6033;
   wire n6034;
   wire n6035;
   wire n6036;
   wire n6037;
   wire n6038;
   wire n6039;
   wire n6040;
   wire n6041;
   wire n6042;
   wire n6043;
   wire n6044;
   wire n6045;
   wire n6046;
   wire n6047;
   wire n6048;
   wire n6049;
   wire n6050;
   wire n6051;
   wire n6052;
   wire n6053;
   wire n6054;
   wire n6055;
   wire n6056;
   wire n6057;
   wire n6058;
   wire n6059;
   wire n6060;
   wire n6061;
   wire n6062;
   wire n6063;
   wire n6064;
   wire n6065;
   wire n6066;
   wire n6067;
   wire n6068;
   wire n6069;
   wire n6070;
   wire n6071;
   wire n6072;
   wire n6073;
   wire n6074;
   wire n6075;
   wire n6076;
   wire n6077;
   wire n6078;
   wire n6079;
   wire n6080;
   wire n6081;
   wire n6082;
   wire n6083;
   wire n6084;
   wire n6085;
   wire n6086;
   wire n6087;
   wire n6088;
   wire n6089;
   wire n6090;
   wire n6091;
   wire n6092;
   wire n6093;
   wire n6094;
   wire n6095;
   wire n6096;
   wire n6097;
   wire n6098;
   wire n6099;
   wire n6100;
   wire n6101;
   wire n6102;
   wire n6103;
   wire n6104;
   wire n6105;
   wire n6106;
   wire n6107;
   wire n6108;
   wire n6109;
   wire n6110;
   wire n6111;
   wire n6112;
   wire n6113;
   wire n6114;
   wire n6115;
   wire n6116;
   wire n6117;
   wire n6118;
   wire n6119;
   wire n6120;
   wire n6121;
   wire n6122;
   wire n6123;
   wire n6124;
   wire n6125;
   wire n6126;
   wire n6127;
   wire n6128;
   wire n6129;
   wire n6130;
   wire n6131;
   wire n6132;
   wire n6133;
   wire n6134;
   wire n6135;
   wire n6136;
   wire n6137;
   wire n6138;
   wire n6139;
   wire n6140;
   wire n6141;
   wire n6142;
   wire n6143;
   wire n6144;
   wire n6145;
   wire n6146;
   wire n6147;
   wire n6148;
   wire n6149;
   wire n6150;
   wire n6151;
   wire n6152;
   wire n6153;
   wire n6154;
   wire n6155;
   wire n6156;
   wire n6157;
   wire n6158;
   wire n6159;
   wire n6160;
   wire n6161;
   wire n6162;
   wire n6163;
   wire n6164;
   wire n6165;
   wire n6166;
   wire n6167;
   wire n6168;
   wire n6169;
   wire n6170;
   wire n6171;
   wire n6172;
   wire n6173;
   wire n6174;
   wire n6175;
   wire n6176;
   wire n6177;
   wire n6178;
   wire n6179;
   wire n6180;
   wire n6181;
   wire n6182;
   wire n6183;
   wire n6184;
   wire n6185;
   wire n6186;
   wire n6187;
   wire n6188;
   wire n6189;
   wire n6190;
   wire n6191;
   wire n6192;
   wire n6193;
   wire n6194;
   wire n6195;
   wire n6196;
   wire n6197;
   wire n6198;
   wire n6199;
   wire n6200;
   wire n6201;
   wire n6202;
   wire n6203;
   wire n6204;
   wire n6205;
   wire n6206;
   wire n6207;
   wire n6208;
   wire n6209;
   wire n6210;
   wire n6211;
   wire n6212;
   wire n6213;
   wire n6214;
   wire n6215;
   wire n6216;
   wire n6217;
   wire n6218;
   wire n6219;
   wire n6220;
   wire n6221;
   wire n6222;
   wire n6223;
   wire n6224;
   wire n6225;
   wire n6226;
   wire n6227;
   wire n6228;
   wire n6229;
   wire n6230;
   wire n6231;
   wire n6232;
   wire n6233;
   wire n6234;
   wire n6235;
   wire n6236;
   wire n6237;
   wire n6238;
   wire n6239;
   wire n6240;
   wire n6241;
   wire n6242;
   wire n6243;
   wire n6244;
   wire n6245;
   wire n6246;
   wire n6247;
   wire n6248;
   wire n6249;
   wire n6250;
   wire n6251;
   wire n6252;
   wire n6253;
   wire n6254;
   wire n6255;
   wire n6256;
   wire n6257;
   wire n6258;
   wire n6259;
   wire n6260;
   wire n6261;
   wire n6262;
   wire n6263;
   wire n6264;
   wire n6265;
   wire n6266;
   wire n6267;
   wire n6268;
   wire n6269;
   wire n6270;
   wire n6271;
   wire n6272;
   wire n6273;
   wire n6274;
   wire n6275;
   wire n6276;
   wire n6277;
   wire n6278;
   wire n6279;
   wire n6280;
   wire n6281;
   wire n6282;
   wire n6283;
   wire n6284;
   wire n6285;
   wire n6286;
   wire n6287;
   wire n6288;
   wire n6289;
   wire n6290;
   wire n6291;
   wire n6292;
   wire n6293;
   wire n6294;
   wire n6295;
   wire n6296;
   wire n6297;
   wire n6298;
   wire n6299;
   wire n6300;
   wire n6301;
   wire n6302;
   wire n6303;
   wire n6304;
   wire n6305;
   wire n6306;
   wire n6307;
   wire n6308;
   wire n6309;
   wire n6310;
   wire n6311;
   wire n6312;
   wire n6313;
   wire n6314;
   wire n6315;
   wire n6316;
   wire n6317;
   wire n6318;
   wire n6319;
   wire n6320;
   wire n6321;
   wire n6322;
   wire n6323;
   wire n6324;
   wire n6325;
   wire n6326;
   wire n6327;
   wire n6328;
   wire n6329;
   wire n6330;
   wire n6331;
   wire n6332;
   wire n6333;
   wire n6334;
   wire n6335;
   wire n6336;
   wire n6337;
   wire n6338;
   wire n6339;
   wire n6340;
   wire n6341;
   wire n6342;
   wire n6343;
   wire n6344;
   wire n6345;
   wire n6346;
   wire n6347;
   wire n6348;
   wire n6349;
   wire n6350;
   wire n6351;
   wire n6352;
   wire n6353;
   wire n6354;
   wire n6355;
   wire n6356;
   wire n6357;
   wire n6358;
   wire n6359;
   wire n6360;
   wire n6361;
   wire n6362;
   wire n6363;
   wire n6364;
   wire n6365;
   wire n6366;
   wire n6367;
   wire n6368;
   wire n6369;
   wire n6370;
   wire n6371;
   wire n6372;
   wire n6373;
   wire n6374;
   wire n6375;
   wire n6376;
   wire n6377;
   wire n6378;
   wire n6379;
   wire n6380;
   wire n6381;
   wire n6382;
   wire n6383;
   wire n6384;
   wire n6385;
   wire n6386;
   wire n6387;
   wire n6388;
   wire n6389;
   wire n6390;
   wire n6391;
   wire n6392;
   wire n6393;
   wire n6394;
   wire n6395;
   wire n6396;
   wire n6397;
   wire n6398;
   wire n6399;
   wire n6400;
   wire n6401;
   wire n6402;
   wire n6403;
   wire n6404;
   wire n6405;
   wire n6406;
   wire n6407;
   wire n6408;
   wire n6409;
   wire n6410;
   wire n6411;
   wire n6412;
   wire n6413;
   wire n6414;
   wire n6415;
   wire n6416;
   wire n6417;
   wire n6418;
   wire n6419;
   wire n6420;
   wire n6421;
   wire n6422;
   wire n6423;
   wire n6424;
   wire n6425;
   wire n6426;
   wire n6427;
   wire n6428;
   wire n6429;
   wire n6430;
   wire n6431;
   wire n6432;
   wire n6433;
   wire n6434;
   wire n6435;
   wire n6436;
   wire n6437;
   wire n6438;
   wire n6439;
   wire n6440;
   wire n6441;
   wire n6442;
   wire n6443;
   wire n6444;
   wire n6445;
   wire n6446;
   wire n6447;
   wire n6448;
   wire n6449;
   wire n6450;
   wire n6451;
   wire n6452;
   wire n6453;
   wire n6454;
   wire n6455;
   wire n6456;
   wire n6457;
   wire n6458;
   wire n6459;
   wire n6460;
   wire n6461;
   wire n6462;
   wire n6463;
   wire n6464;
   wire n6465;
   wire n6466;
   wire n6467;
   wire n6468;
   wire n6469;
   wire n6470;
   wire n6471;
   wire n6472;
   wire n6473;
   wire n6474;
   wire n6475;
   wire n6476;
   wire n6477;
   wire n6478;
   wire n6479;
   wire n6480;
   wire n6481;
   wire n6482;
   wire n6483;
   wire n6484;
   wire n6485;
   wire n6486;
   wire n6487;
   wire n6488;
   wire n6489;
   wire n6490;
   wire n6491;
   wire n6492;
   wire n6493;
   wire n6494;
   wire n6495;
   wire n6496;
   wire n6497;
   wire n6498;
   wire n6499;
   wire n6500;
   wire n6501;
   wire n6502;
   wire n6503;
   wire n6504;
   wire n6505;
   wire n6506;
   wire n6507;
   wire n6508;
   wire n6509;
   wire n6510;
   wire n6511;
   wire n6512;
   wire n6513;
   wire n6514;
   wire n6515;
   wire n6516;
   wire n6517;
   wire n6518;
   wire n6519;
   wire n6520;
   wire n6521;
   wire n6522;
   wire n6523;
   wire n6524;
   wire n6525;
   wire n6526;
   wire n6527;
   wire n6528;
   wire n6529;
   wire n6530;
   wire n6531;
   wire n6532;
   wire n6533;
   wire n6534;
   wire n6535;
   wire n6536;
   wire n6537;
   wire n6538;
   wire n6539;
   wire n6540;
   wire n6541;
   wire n6542;
   wire n6543;
   wire n6544;
   wire n6545;
   wire n6546;
   wire n6547;
   wire n6548;
   wire n6549;
   wire n6550;
   wire n6551;
   wire n6552;
   wire n6553;
   wire n6554;
   wire n6555;
   wire n6556;
   wire n6557;
   wire n6558;
   wire n6559;
   wire n6560;
   wire n6561;
   wire n6562;
   wire n6563;
   wire n6564;
   wire n6565;
   wire n6566;
   wire n6567;
   wire n6568;
   wire n6569;
   wire n6570;
   wire n6571;
   wire n6572;
   wire n6573;
   wire n6574;
   wire n6575;
   wire n6576;
   wire n6577;
   wire n6578;
   wire n6579;
   wire n6580;
   wire n6581;
   wire n6582;
   wire n6583;
   wire n6584;
   wire n6585;
   wire n6586;
   wire n6587;
   wire n6588;
   wire n6589;
   wire n6590;
   wire n6591;
   wire n6592;
   wire n6593;
   wire n6594;
   wire n6595;
   wire n6596;
   wire n6597;
   wire n6598;
   wire n6599;
   wire n6600;
   wire n6601;
   wire n6602;
   wire n6603;
   wire n6604;
   wire n6605;
   wire n6606;
   wire n6607;
   wire n6608;
   wire n6609;
   wire n6610;
   wire n6611;
   wire n6612;
   wire n6613;
   wire n6614;
   wire n6615;
   wire n6616;
   wire n6617;
   wire n6618;
   wire n6619;
   wire n6620;
   wire n6621;
   wire n6622;
   wire n6623;
   wire n6624;
   wire n6625;
   wire n6626;
   wire n6627;
   wire n6628;
   wire n6629;
   wire n6630;
   wire n6631;
   wire n6632;
   wire n6633;
   wire n6634;
   wire n6635;
   wire n6636;
   wire n6637;
   wire n6638;
   wire n6639;
   wire n6640;
   wire n6641;
   wire n6642;
   wire n6643;
   wire n6644;
   wire n6645;
   wire n6646;
   wire n6647;
   wire n6648;
   wire n6649;
   wire n6650;
   wire n6651;
   wire n6652;
   wire n6653;
   wire n6654;
   wire n6655;
   wire n6656;
   wire n6657;
   wire n6658;
   wire n6659;
   wire n6660;
   wire n6661;
   wire n6662;
   wire n6663;
   wire n6664;
   wire n6665;
   wire n6666;
   wire n6667;
   wire n6668;
   wire n6669;
   wire n6670;
   wire n6671;
   wire n6672;
   wire n6673;
   wire n6674;
   wire n6675;
   wire n6676;
   wire n6677;
   wire n6678;
   wire n6679;
   wire n6680;
   wire n6681;
   wire n6682;
   wire n6683;
   wire n6684;
   wire n6685;
   wire n6686;
   wire n6687;
   wire n6688;
   wire n6689;
   wire n6690;
   wire n6691;
   wire n6692;
   wire n6693;
   wire n6694;
   wire n6695;
   wire n6696;
   wire n6697;
   wire n6698;
   wire n6699;
   wire n6700;
   wire n6701;
   wire n6702;
   wire n6703;
   wire n6704;
   wire n6705;
   wire n6706;
   wire n6707;
   wire n6708;
   wire n6709;
   wire n6710;
   wire n6711;
   wire n6712;
   wire n6713;
   wire n6714;
   wire n6715;
   wire n6716;
   wire n6717;
   wire n6718;
   wire n6719;
   wire n6720;
   wire n6721;
   wire n6722;
   wire n6723;
   wire n6724;
   wire n6725;
   wire n6726;
   wire n6727;
   wire n6728;
   wire n6729;
   wire n6730;
   wire n6731;
   wire n6732;
   wire n6733;
   wire n6734;
   wire n6735;
   wire n6736;
   wire n6737;
   wire n6738;
   wire n6739;
   wire n6740;
   wire n6741;
   wire n6742;
   wire n6743;
   wire n6744;
   wire n6745;
   wire n6746;
   wire n6747;
   wire n6748;
   wire n6749;
   wire n6750;
   wire n6751;
   wire n6752;
   wire n6753;
   wire n6754;
   wire n6755;
   wire n6756;
   wire n6757;
   wire n6758;
   wire n6759;
   wire n6760;
   wire n6761;
   wire n6762;
   wire n6763;
   wire n6764;
   wire n6765;
   wire n6766;
   wire \add_x_22_5/carry[2] ;
   wire \add_x_22_5/carry[3] ;
   wire \add_x_22_5/carry[4] ;
   wire \add_x_22_5/carry[5] ;
   wire \add_x_22_5/carry[6] ;
   wire \add_x_22_5/carry[7] ;
   wire \add_x_22_5/carry[8] ;
   wire \add_x_22_5/carry[9] ;
   wire \add_x_22_5/carry[10] ;
   wire \add_x_22_5/carry[11] ;
   wire \add_x_22_5/carry[12] ;
   wire \add_x_22_5/carry[13] ;
   wire \add_x_22_5/carry[14] ;
   wire \add_x_22_5/carry[15] ;
   wire \add_x_22_5/carry[16] ;
   wire \add_x_22_5/carry[17] ;
   wire \add_x_22_5/carry[18] ;
   wire \add_x_22_5/carry[19] ;
   wire \add_x_22_5/carry[20] ;
   wire \add_x_22_5/carry[21] ;
   wire \add_x_22_5/carry[22] ;
   wire \add_x_22_5/carry[23] ;
   wire \add_x_22_5/carry[24] ;
   wire \add_x_22_5/carry[25] ;
   wire \add_x_22_5/carry[26] ;
   wire \add_x_22_5/carry[27] ;
   wire \add_x_22_5/carry[28] ;
   wire \add_x_22_5/carry[29] ;
   wire \add_x_22_5/carry[30] ;
   wire \add_x_22_5/carry[31] ;
   wire \add_x_22_3/carry[2] ;
   wire \add_x_22_3/carry[3] ;
   wire \add_x_22_3/carry[4] ;
   wire \add_x_22_3/carry[5] ;
   wire \add_x_22_3/carry[6] ;
   wire \add_x_22_3/carry[7] ;
   wire \add_x_22_3/carry[8] ;
   wire \add_x_22_3/carry[9] ;
   wire \add_x_22_3/carry[10] ;
   wire \add_x_22_3/carry[11] ;
   wire \add_x_22_3/carry[12] ;
   wire \add_x_22_3/carry[13] ;
   wire \add_x_22_3/carry[14] ;
   wire \add_x_22_3/carry[15] ;
   wire \add_x_22_3/carry[16] ;
   wire \add_x_22_3/carry[17] ;
   wire \add_x_22_3/carry[18] ;
   wire \add_x_22_3/carry[19] ;
   wire \add_x_22_3/carry[20] ;
   wire \add_x_22_3/carry[21] ;
   wire \add_x_22_3/carry[22] ;
   wire \add_x_22_3/carry[23] ;
   wire \add_x_22_3/carry[24] ;
   wire \add_x_22_3/carry[25] ;
   wire \add_x_22_3/carry[26] ;
   wire \add_x_22_3/carry[27] ;
   wire \add_x_22_3/carry[28] ;
   wire \add_x_22_3/carry[29] ;
   wire \add_x_22_3/carry[30] ;
   wire \add_x_22_3/carry[31] ;
   wire \add_x_22_2/carry[2] ;
   wire \add_x_22_2/carry[3] ;
   wire \add_x_22_2/carry[4] ;
   wire \add_x_22_2/carry[5] ;
   wire \add_x_22_2/carry[6] ;
   wire \add_x_22_2/carry[7] ;
   wire \add_x_22_2/carry[8] ;
   wire \add_x_22_2/carry[9] ;
   wire \add_x_22_2/carry[10] ;
   wire \add_x_22_2/carry[11] ;
   wire \add_x_22_2/carry[12] ;
   wire \add_x_22_2/carry[13] ;
   wire \add_x_22_2/carry[14] ;
   wire \add_x_22_2/carry[15] ;
   wire \add_x_22_2/carry[16] ;
   wire \add_x_22_2/carry[17] ;
   wire \add_x_22_2/carry[18] ;
   wire \add_x_22_2/carry[19] ;
   wire \add_x_22_2/carry[20] ;
   wire \add_x_22_2/carry[21] ;
   wire \add_x_22_2/carry[22] ;
   wire \add_x_22_2/carry[23] ;
   wire \add_x_22_2/carry[24] ;
   wire \add_x_22_2/carry[25] ;
   wire \add_x_22_2/carry[26] ;
   wire \add_x_22_2/carry[27] ;
   wire \add_x_22_2/carry[28] ;
   wire \add_x_22_2/carry[29] ;
   wire \add_x_22_2/carry[30] ;
   wire \add_x_22_2/carry[31] ;
   wire \add_x_22_1/carry[2] ;
   wire \add_x_22_1/carry[3] ;
   wire \add_x_22_1/carry[4] ;
   wire \add_x_22_1/carry[5] ;
   wire \add_x_22_1/carry[6] ;
   wire \add_x_22_1/carry[7] ;
   wire \add_x_22_1/carry[8] ;
   wire \add_x_22_1/carry[9] ;
   wire \add_x_22_1/carry[10] ;
   wire \add_x_22_1/carry[11] ;
   wire \add_x_22_1/carry[12] ;
   wire \add_x_22_1/carry[13] ;
   wire \add_x_22_1/carry[14] ;
   wire \add_x_22_1/carry[15] ;
   wire \add_x_22_1/carry[16] ;
   wire \add_x_22_1/carry[17] ;
   wire \add_x_22_1/carry[18] ;
   wire \add_x_22_1/carry[19] ;
   wire \add_x_22_1/carry[20] ;
   wire \add_x_22_1/carry[21] ;
   wire \add_x_22_1/carry[22] ;
   wire \add_x_22_1/carry[23] ;
   wire \add_x_22_1/carry[24] ;
   wire \add_x_22_1/carry[25] ;
   wire \add_x_22_1/carry[26] ;
   wire \add_x_22_1/carry[27] ;
   wire \add_x_22_1/carry[28] ;
   wire \add_x_22_1/carry[29] ;
   wire \add_x_22_1/carry[30] ;
   wire \add_x_22_1/carry[31] ;
   wire \add_x_22_0/carry[2] ;
   wire \add_x_22_0/carry[3] ;
   wire \add_x_22_0/carry[4] ;
   wire \add_x_22_0/carry[5] ;
   wire \add_x_22_0/carry[6] ;
   wire \add_x_22_0/carry[7] ;
   wire \add_x_22_0/carry[8] ;
   wire \add_x_22_0/carry[9] ;
   wire \add_x_22_0/carry[10] ;
   wire \add_x_22_0/carry[11] ;
   wire \add_x_22_0/carry[12] ;
   wire \add_x_22_0/carry[13] ;
   wire \add_x_22_0/carry[14] ;
   wire \add_x_22_0/carry[15] ;
   wire \add_x_22_0/carry[16] ;
   wire \add_x_22_0/carry[17] ;
   wire \add_x_22_0/carry[18] ;
   wire \add_x_22_0/carry[19] ;
   wire \add_x_22_0/carry[20] ;
   wire \add_x_22_0/carry[21] ;
   wire \add_x_22_0/carry[22] ;
   wire \add_x_22_0/carry[23] ;
   wire \add_x_22_0/carry[24] ;
   wire \add_x_22_0/carry[25] ;
   wire \add_x_22_0/carry[26] ;
   wire \add_x_22_0/carry[27] ;
   wire \add_x_22_0/carry[28] ;
   wire \add_x_22_0/carry[29] ;
   wire \add_x_22_0/carry[30] ;
   wire \add_x_22_0/carry[31] ;
   wire n6768;
   wire n6769;
   wire n6770;
   wire n6771;
   wire n6772;
   wire n6773;
   wire n6774;
   wire n6775;
   wire n6776;
   wire n6777;
   wire n6778;
   wire n6779;
   wire n6780;
   wire n6781;
   wire n6782;
   wire n6783;
   wire n6784;
   wire n6785;
   wire n6786;
   wire n6787;
   wire n6788;
   wire n6789;
   wire n6790;
   wire n6791;
   wire n6792;
   wire n6793;
   wire n6794;
   wire n6795;
   wire n6796;
   wire n6797;
   wire n6798;
   wire n6799;
   wire n6800;
   wire n6801;
   wire n6802;
   wire n6803;
   wire n6804;
   wire n6805;
   wire n6806;
   wire n6807;
   wire n6808;
   wire n6809;
   wire n6810;
   wire n6811;
   wire n6812;
   wire n6813;
   wire n6814;
   wire n6815;
   wire n6816;
   wire n6817;
   wire n6818;
   wire n6819;
   wire n6820;
   wire n6821;
   wire n6822;
   wire n6823;
   wire n6824;
   wire n6825;
   wire n6826;
   wire n6827;
   wire n6828;
   wire n6829;
   wire n6830;
   wire n6831;
   wire n6832;
   wire n6833;
   wire n6834;
   wire n6835;
   wire n6836;
   wire n6837;
   wire n6838;
   wire n6839;
   wire n6840;
   wire n6841;
   wire n6842;
   wire n6843;
   wire n6844;
   wire n6845;
   wire n6846;
   wire n6847;
   wire n6848;
   wire n6849;
   wire n6850;
   wire n6851;
   wire n6852;
   wire n6853;
   wire n6854;
   wire n6855;
   wire n6856;
   wire n6857;
   wire n6858;
   wire n6859;
   wire n6860;
   wire n6861;
   wire n6862;
   wire n6863;
   wire n6864;
   wire n6865;
   wire n6866;
   wire n6867;
   wire n6868;
   wire n6869;
   wire n6870;
   wire n6871;
   wire n6872;
   wire n6873;
   wire n6874;
   wire n6875;
   wire n6876;
   wire n6877;
   wire n6878;
   wire n6879;
   wire n6880;
   wire n6881;
   wire n6882;
   wire n6883;
   wire n6884;
   wire n6885;
   wire n6886;
   wire n6887;
   wire n6888;
   wire n6889;
   wire n6890;
   wire n6891;
   wire n6892;
   wire n6893;
   wire n6894;
   wire n6895;
   wire n6896;
   wire n6897;
   wire n6898;
   wire n6899;
   wire n6900;
   wire n6901;
   wire n6902;
   wire n6903;
   wire n6904;
   wire n6905;
   wire n6906;
   wire n6907;
   wire n6908;
   wire n6909;
   wire n6910;
   wire n6911;
   wire n6912;
   wire n6913;
   wire n6914;
   wire n6915;
   wire n6916;
   wire n6917;
   wire n6918;
   wire n6919;
   wire n6920;
   wire n6921;
   wire n6922;
   wire n6923;
   wire n6924;
   wire n6925;
   wire n6926;
   wire n6927;
   wire n6928;
   wire n6929;
   wire n6930;
   wire n6931;
   wire n6932;
   wire n6933;
   wire n6934;
   wire n6935;
   wire n6936;
   wire n6937;
   wire n6938;
   wire n6939;
   wire n6940;
   wire n6941;
   wire n6942;
   wire n6943;
   wire n6944;
   wire n6945;
   wire n6946;
   wire n6947;
   wire n6948;
   wire n6949;
   wire n6950;
   wire n6951;
   wire n6952;
   wire n6953;
   wire n6954;
   wire n6955;
   wire n6956;
   wire n6957;
   wire n6958;
   wire n6959;
   wire n6960;
   wire n6961;
   wire n6962;
   wire n6963;
   wire n6964;
   wire n6965;
   wire n6966;
   wire n6967;
   wire n6968;
   wire n6969;
   wire n6970;
   wire n6971;
   wire n6972;
   wire n6973;
   wire n6974;
   wire n6975;
   wire n6976;
   wire n6977;
   wire n6978;
   wire n6979;
   wire n6980;
   wire n6981;
   wire n6982;
   wire n6983;
   wire n6984;
   wire n6985;
   wire n6986;
   wire n6987;
   wire n6988;
   wire n6989;
   wire n6990;
   wire n6991;
   wire n6992;
   wire n6993;
   wire n6994;
   wire n6995;
   wire n6996;
   wire n6997;
   wire n6998;
   wire n6999;
   wire n7000;
   wire n7001;
   wire n7002;
   wire n7003;
   wire n7004;
   wire n7005;
   wire n7006;
   wire n7007;
   wire n7008;
   wire n7009;
   wire n7010;
   wire n7011;
   wire n7012;
   wire n7013;
   wire n7014;
   wire n7015;
   wire n7016;
   wire n7017;
   wire n7018;
   wire n7019;
   wire n7020;
   wire n7021;
   wire n7022;
   wire n7023;
   wire n7056;
   wire n7057;
   wire n7058;
   wire n7059;
   wire n7060;
   wire n7061;
   wire n7062;
   wire n7063;
   wire n7064;
   wire n7065;
   wire n7066;
   wire n7067;
   wire n7068;
   wire n7069;
   wire n7070;
   wire n7071;
   wire n7072;
   wire n7073;
   wire n7074;
   wire n7075;
   wire n7076;
   wire n7077;
   wire n7078;
   wire n7079;
   wire n7080;
   wire n7081;
   wire n7082;
   wire n7083;
   wire n7084;
   wire n7085;
   wire n7086;
   wire n7087;
   wire n7088;
   wire n7089;
   wire n7090;
   wire n7091;
   wire n7092;
   wire n7093;
   wire n7094;
   wire n7095;
   wire n7096;
   wire n7097;
   wire n7098;
   wire n7099;
   wire n7100;
   wire n7101;
   wire n7102;
   wire n7103;
   wire n7104;
   wire n7105;
   wire n7106;
   wire n7107;
   wire n7108;
   wire n7109;
   wire n7110;
   wire n7111;
   wire n7112;
   wire n7113;
   wire n7114;
   wire n7115;
   wire n7116;
   wire n7117;
   wire n7118;
   wire n7119;
   wire n7120;
   wire n7121;
   wire n7122;
   wire n7123;
   wire n7124;
   wire n7125;
   wire n7126;
   wire n7127;
   wire n7128;
   wire n7129;
   wire n7130;
   wire n7131;
   wire n7132;
   wire n7133;
   wire n7134;
   wire n7135;
   wire n7136;
   wire n7137;
   wire n7138;
   wire n7139;
   wire n7140;
   wire n7141;
   wire n7142;
   wire n7143;
   wire n7144;
   wire n7145;
   wire n7146;
   wire n7147;
   wire n7148;
   wire n7149;
   wire n7150;
   wire n7151;
   wire n7152;
   wire n7153;
   wire n7154;
   wire n7155;
   wire n7156;
   wire n7157;
   wire n7158;
   wire n7159;
   wire n7160;
   wire n7161;
   wire n7162;
   wire n7163;
   wire n7164;
   wire n7165;
   wire n7166;
   wire n7167;
   wire n7168;
   wire n7169;
   wire n7170;
   wire n7171;
   wire n7172;
   wire n7173;
   wire n7174;
   wire n7175;
   wire n7176;
   wire n7177;
   wire n7178;
   wire n7179;
   wire n7180;
   wire n7181;
   wire n7182;
   wire n7183;
   wire n7184;
   wire n7185;
   wire n7186;
   wire n7187;
   wire n7188;
   wire n7189;
   wire n7190;
   wire n7191;
   wire n7192;
   wire n7193;
   wire n7194;
   wire n7195;
   wire n7196;
   wire n7197;
   wire n7198;
   wire n7199;
   wire n7200;
   wire n7201;
   wire n7202;
   wire n7203;
   wire n7204;
   wire n7205;
   wire n7206;
   wire n7207;
   wire n7208;
   wire n7209;
   wire n7210;
   wire n7211;
   wire n7212;
   wire n7213;
   wire n7214;
   wire n7215;
   wire n7216;
   wire n7217;
   wire n7218;
   wire n7219;
   wire n7220;
   wire n7221;
   wire n7222;
   wire n7223;
   wire n7224;
   wire n7225;
   wire n7226;
   wire n7227;
   wire n7228;
   wire n7229;
   wire n7230;
   wire n7231;
   wire n7232;
   wire n7233;
   wire n7234;
   wire n7235;
   wire n7236;
   wire n7237;
   wire n7238;
   wire n7239;
   wire n7240;
   wire n7241;
   wire n7242;
   wire n7243;
   wire n7244;
   wire n7245;
   wire n7246;
   wire n7247;
   wire n7248;
   wire n7249;
   wire n7250;
   wire n7251;
   wire n7252;
   wire n7253;
   wire n7254;
   wire n7255;
   wire n7256;
   wire n7257;
   wire n7258;
   wire n7259;
   wire n7260;
   wire n7261;
   wire n7262;
   wire n7263;
   wire n7264;
   wire n7265;
   wire n7266;
   wire n7267;
   wire n7268;
   wire n7269;
   wire n7270;
   wire n7271;
   wire n7272;
   wire n7273;
   wire n7274;
   wire n7275;
   wire n7276;
   wire n7277;
   wire n7278;
   wire n7279;
   wire n7280;
   wire n7281;
   wire n7282;
   wire n7283;
   wire n7284;
   wire n7285;
   wire n7286;
   wire n7287;
   wire n7288;
   wire n7289;
   wire n7290;
   wire n7291;
   wire n7292;
   wire n7293;
   wire n7294;
   wire n7295;
   wire n7297;
   wire n7298;
   wire n7299;
   wire n7300;
   wire n7301;
   wire n7302;
   wire n7303;
   wire n7304;
   wire n7305;
   wire n7306;
   wire n7307;
   wire n7308;
   wire n7309;
   wire n7310;
   wire n7311;
   wire n7312;
   wire n7313;
   wire n7314;
   wire n7315;
   wire n7316;
   wire n7317;
   wire n7318;
   wire n7319;
   wire n7320;
   wire n7321;
   wire n7322;
   wire n7323;
   wire n7324;
   wire n7325;
   wire n7326;
   wire n7327;
   wire n7328;
   wire n7329;
   wire n7330;
   wire n7331;
   wire n7332;
   wire n7333;
   wire n7334;
   wire n7335;
   wire n7336;
   wire n7337;
   wire n7338;
   wire n7339;
   wire n7340;
   wire n7341;
   wire n7342;
   wire n7343;
   wire n7344;
   wire n7345;
   wire n7346;
   wire n7347;
   wire n7348;
   wire n7349;
   wire n7350;
   wire n7351;
   wire n7352;
   wire n7353;
   wire n7354;
   wire n7355;
   wire n7356;
   wire n7357;
   wire n7358;
   wire n7359;
   wire n7360;
   wire n7361;
   wire n7362;
   wire n7363;
   wire n7364;
   wire n7365;
   wire n7366;
   wire n7367;
   wire n7368;
   wire n7369;
   wire n7370;
   wire n7371;
   wire n7372;
   wire n7373;
   wire n7374;
   wire n7375;
   wire n7376;
   wire n7377;
   wire n7378;
   wire n7379;
   wire n7380;
   wire n7381;
   wire n7382;
   wire n7383;
   wire n7384;
   wire n7385;
   wire n7386;
   wire n7387;
   wire n7388;
   wire n7389;
   wire n7390;
   wire n7391;
   wire n7392;
   wire n7393;
   wire n7394;
   wire n7395;
   wire n7396;
   wire n7397;
   wire n7398;
   wire n7399;
   wire n7400;
   wire n7401;
   wire n7402;
   wire n7403;
   wire n7404;
   wire n7405;
   wire n7406;
   wire n7407;
   wire n7408;
   wire n7409;
   wire n7410;
   wire n7411;
   wire n7412;
   wire n7413;
   wire n7414;
   wire n7415;
   wire n7416;
   wire n7417;
   wire n7418;
   wire n7419;
   wire n7420;
   wire n7421;
   wire n7422;
   wire n7423;
   wire n7424;
   wire n7425;
   wire n7426;
   wire n7427;
   wire n7428;
   wire n7429;
   wire n7430;
   wire n7431;
   wire n7432;
   wire n7433;
   wire n7434;
   wire n7435;
   wire n7436;
   wire n7437;
   wire n7438;
   wire n7439;
   wire n7440;
   wire n7441;
   wire n7442;
   wire n7443;
   wire n7444;
   wire n7445;
   wire n7446;
   wire n7447;
   wire n7448;
   wire n7449;
   wire n7450;
   wire n7451;
   wire n7452;
   wire n7453;
   wire n7454;
   wire n7455;
   wire n7456;
   wire n7457;
   wire n7458;
   wire n7459;
   wire n7460;
   wire n7461;
   wire n7462;
   wire n7463;
   wire n7464;
   wire n7465;
   wire n7466;
   wire n7467;
   wire n7468;
   wire n7469;
   wire n7470;
   wire n7471;
   wire n7472;
   wire n7473;
   wire n7474;
   wire n7475;
   wire n7476;
   wire n7477;
   wire n7478;
   wire n7479;
   wire n7480;
   wire n7481;
   wire n7482;
   wire n7483;
   wire n7484;
   wire n7485;
   wire n7486;
   wire n7487;
   wire n7488;
   wire n7489;
   wire n7490;
   wire n7491;
   wire n7492;
   wire n7493;
   wire n7494;
   wire n7495;
   wire n7496;
   wire n7497;
   wire n7498;
   wire n7499;
   wire n7500;
   wire n7501;
   wire n7502;
   wire n7503;
   wire n7504;
   wire n7505;
   wire n7506;
   wire n7507;
   wire n7508;
   wire n7509;
   wire n7510;
   wire n7511;
   wire n7512;
   wire n7513;
   wire n7514;
   wire n7515;
   wire n7516;
   wire n7517;
   wire n7518;
   wire n7519;
   wire n7520;
   wire n7521;
   wire n7522;
   wire n7523;
   wire n7524;
   wire n7525;
   wire n7526;
   wire n7527;
   wire n7528;
   wire n7529;
   wire n7530;
   wire n7531;
   wire n7532;
   wire n7533;
   wire n7534;
   wire n7535;
   wire n7536;
   wire n7537;
   wire n7538;
   wire n7539;
   wire n7540;
   wire n7541;
   wire n7542;
   wire n7543;
   wire n7544;
   wire n7545;
   wire n7546;
   wire n7547;
   wire n7548;
   wire n7549;
   wire n7550;
   wire n7551;
   wire n7552;
   wire n7553;
   wire n7554;
   wire n7555;
   wire n7556;
   wire n7557;
   wire n7558;
   wire n7559;
   wire n7560;
   wire n7561;
   wire n7562;
   wire n7563;
   wire n7564;
   wire n7565;
   wire n7566;
   wire n7567;
   wire n7568;
   wire n7569;
   wire n7570;
   wire n7571;
   wire n7572;
   wire n7573;
   wire n7574;
   wire n7575;
   wire n7576;
   wire n7577;
   wire n7578;
   wire n7579;
   wire n7580;
   wire n7581;
   wire n7582;
   wire n7583;
   wire n7584;
   wire n7585;
   wire n7586;
   wire n7587;
   wire n7588;
   wire n7589;
   wire n7590;
   wire n7591;
   wire n7592;
   wire n7593;
   wire n7594;
   wire n7595;
   wire n7596;
   wire n7597;
   wire n7598;
   wire n7599;
   wire n7600;
   wire n7601;
   wire n7602;
   wire n7603;
   wire n7606;
   wire n7607;
   wire n7608;
   wire n7609;
   wire n7610;
   wire n7611;
   wire n7614;
   wire n7615;
   wire n7616;
   wire n7617;
   wire n7618;
   wire n7619;
   wire n7952;
   wire n7953;
   wire n7955;
   wire n7956;
   wire n7957;
   wire n7958;
   wire n7959;
   wire n7960;
   wire n7962;
   wire n7963;
   wire n7964;
   wire n7965;
   wire n7966;
   wire n7967;
   wire n7968;
   wire n7969;
   wire n7970;
   wire n7971;
   wire n7972;
   wire n7973;
   wire n7974;
   wire n7975;
   wire n7976;
   wire n7977;
   wire n8011;
   wire n8012;
   wire n8013;
   wire n8014;
   wire n8015;
   wire n8016;
   wire n8017;
   wire n8018;
   wire n8019;
   wire n8020;
   wire n8021;
   wire n8022;
   wire n8023;
   wire n8024;
   wire n8025;
   wire n8026;
   wire n8027;
   wire n8028;
   wire n8029;
   wire n8030;
   wire n8031;
   wire n8032;
   wire n8033;
   wire n8034;
   wire n8035;
   wire n8036;
   wire n8037;
   wire n8038;
   wire n8039;
   wire n8040;
   wire n8041;
   wire n8042;
   wire n8050;
   wire n8051;
   wire n8052;
   wire n8053;
   wire n8054;
   wire n8055;
   wire n8056;
   wire n8057;
   wire n8058;
   wire n8059;
   wire n8060;
   wire n8061;
   wire n8062;
   wire n8063;
   wire n8064;
   wire n8065;
   wire n8066;
   wire n8067;
   wire n8068;
   wire n8069;
   wire n8070;
   wire n8071;
   wire n8072;
   wire n8073;
   wire n8074;
   wire n8075;
   wire n8076;
   wire n8077;
   wire n8078;
   wire n8079;
   wire n8080;
   wire n8081;
   wire n8082;
   wire n8083;
   wire n8084;
   wire n8085;
   wire n8086;
   wire n8087;
   wire n8088;
   wire n8089;
   wire n8090;
   wire n8091;
   wire n8092;
   wire n8093;
   wire n8094;
   wire n8095;
   wire n8137;
   wire n8138;
   wire n8139;
   wire n8140;
   wire n8141;
   wire n8142;
   wire n8143;
   wire n8144;
   wire n8145;
   wire n8376;
   wire n8377;
   wire n8378;
   wire n8379;
   wire n8380;
   wire n8381;
   wire n8382;
   wire n8383;
   wire n8384;
   wire n8472;
   wire n8473;
   wire n8474;
   wire n8475;
   wire n8476;
   wire n8477;
   wire n8478;
   wire n8479;
   wire n8480;
   wire n8711;
   wire n8712;
   wire n8713;
   wire n8714;
   wire n8715;
   wire n8716;
   wire n8717;
   wire n8718;
   wire n8719;
   wire n8784;
   wire n8785;
   wire n8786;
   wire n8787;
   wire n8788;
   wire n8789;
   wire n8790;
   wire n8791;
   wire n8805;
   wire n8806;
   wire n8807;
   wire n8808;
   wire n8809;
   wire n8810;
   wire n8811;
   wire n8812;
   wire n8837;
   wire n8838;
   wire n8839;
   wire n8840;
   wire n8841;
   wire n8842;
   wire n8843;
   wire n8844;
   wire n8845;
   wire n8870;
   wire n8871;
   wire n8872;
   wire n8873;
   wire n8874;
   wire n8875;
   wire n8876;
   wire n8877;
   wire n8878;
   wire n9370;
   wire n9371;
   wire n9372;
   wire n9373;
   wire n9374;
   wire n9375;
   wire n9376;
   wire n9377;
   wire n9378;
   wire n9381;
   wire n9382;
   wire n9383;
   wire n9384;
   wire n9385;
   wire n9386;
   wire n9387;
   wire n9388;
   wire n9389;
   wire n9390;
   wire n9391;
   wire n9406;
   wire n9407;
   wire n9408;
   wire n9409;
   wire n9410;
   wire n9411;
   wire n9412;
   wire n9413;
   wire n9414;
   wire n9415;
   wire n9416;
   wire n9417;
   wire n9418;
   wire n9419;
   wire n9420;
   wire n9421;
   wire n9431;
   wire n9432;
   wire n9433;
   wire n9434;
   wire n9435;
   wire n9436;
   wire n9437;
   wire n9438;
   wire n9439;
   wire n9440;
   wire n9441;
   wire n9442;
   wire n9443;
   wire n9444;
   wire n9445;
   wire n9446;
   wire n9447;
   wire n9448;
   wire n9449;
   wire n9462;
   wire n9463;
   wire n9464;
   wire n9465;
   wire n9466;
   wire n9467;
   wire n9468;
   wire n9469;
   wire n9470;
   wire n9471;
   wire n9472;
   wire n9473;
   wire n9474;
   wire n9475;
   wire n9476;
   wire n9477;
   wire n9478;
   wire n9479;
   wire n9480;
   wire n9481;
   wire n9482;
   wire n9483;
   wire n9484;
   wire n9485;
   wire n9486;
   wire n9487;
   wire n9488;
   wire n9489;
   wire n9490;
   wire n9491;
   wire n9492;
   wire n9493;
   wire n9494;
   wire n9495;
   wire n9496;
   wire n9497;
   wire n9498;
   wire n9499;
   wire n9500;
   wire n9501;
   wire n9502;
   wire n9503;
   wire n9504;
   wire n9505;
   wire n9506;
   wire n9507;
   wire n9508;
   wire n9509;
   wire n9510;
   wire n9511;
   wire n9512;
   wire n9513;
   wire n9514;
   wire n9515;
   wire n9516;
   wire n9517;
   wire n9518;
   wire n9519;
   wire n9520;
   wire n9521;
   wire n9522;
   wire n9523;
   wire n9524;
   wire n9525;
   wire n9526;
   wire n9527;
   wire n9528;
   wire n9529;
   wire n9530;
   wire n9531;
   wire n9532;
   wire n9533;
   wire n9534;
   wire n9535;
   wire n9536;
   wire n9537;
   wire n9538;
   wire n9539;
   wire n9540;
   wire n9541;
   wire n9542;
   wire n9543;
   wire n9544;
   wire n9545;
   wire n9546;
   wire n9547;
   wire [31:0] instruction;
   wire [31:0] fft_data_in;
   wire [31:0] fir_data_in;

   CLKINVX16TS clk__L1_I0 (.Y(clk__L1_N0), 
	.A(clk));
   CLKBUFX2TS FE_OFC1825_n7107 (.Y(FE_OFN1825_n7107), 
	.A(n7107));
   CLKBUFX2TS FE_OFC1824_router_addr_calc_fir_read_calc_count_5_ (.Y(FE_OFN1824_router_addr_calc_fir_read_calc_count_5_), 
	.A(\router/addr_calc/fir_read_calc/count[5] ));
   CLKBUFX2TS FE_OFC1823_n4643 (.Y(FE_OFN1823_n4643), 
	.A(FE_OFN719_n4643));
   CLKBUFX2TS FE_OFC1822_n4643 (.Y(FE_OFN1822_n4643), 
	.A(FE_OFN721_n4643));
   CLKINVX1TS FE_OFC1821_acc_fft_data_in_28_ (.Y(FE_OFN1821_acc_fft_data_in_28_), 
	.A(FE_OFN1819_acc_fft_data_in_28_));
   CLKINVX1TS FE_OFC1820_acc_fft_data_in_28_ (.Y(FE_OFN1820_acc_fft_data_in_28_), 
	.A(FE_OFN1819_acc_fft_data_in_28_));
   CLKINVX1TS FE_OFC1819_acc_fft_data_in_28_ (.Y(FE_OFN1819_acc_fft_data_in_28_), 
	.A(FE_OFN1469_acc_fft_data_in_28_));
   CLKBUFX2TS FE_OFC1818_acc_fir_data_in_26_ (.Y(FE_OFN1818_acc_fir_data_in_26_), 
	.A(FE_OFN1656_acc_fir_data_in_26_));
   BUFX2TS FE_MDBC15_U5584 (.Y(FE_MDBN15_), 
	.A(fft_data_in[7]));
   CLKINVX1TS FE_OFC1817_acc_fir_data_in_0_ (.Y(FE_OFN1817_acc_fir_data_in_0_), 
	.A(FE_OFN1815_acc_fir_data_in_0_));
   CLKINVX1TS FE_OFC1816_acc_fir_data_in_0_ (.Y(FE_OFN1816_acc_fir_data_in_0_), 
	.A(FE_OFN1815_acc_fir_data_in_0_));
   CLKINVX1TS FE_OFC1815_acc_fir_data_in_0_ (.Y(FE_OFN1815_acc_fir_data_in_0_), 
	.A(FE_OFN1813_acc_fir_data_in_0_));
   CLKBUFX2TS FE_OFC1814_acc_fir_data_in_0_ (.Y(FE_OFN1814_acc_fir_data_in_0_), 
	.A(FE_OFN1811_acc_fir_data_in_0_));
   CLKBUFX2TS FE_OFC1813_acc_fir_data_in_0_ (.Y(FE_OFN1813_acc_fir_data_in_0_), 
	.A(FE_OFN1811_acc_fir_data_in_0_));
   CLKINVX1TS FE_OFC1812_acc_fir_data_in_0_ (.Y(FE_OFN1812_acc_fir_data_in_0_), 
	.A(FE_OFN1809_acc_fir_data_in_0_));
   CLKINVX1TS FE_OFC1811_acc_fir_data_in_0_ (.Y(FE_OFN1811_acc_fir_data_in_0_), 
	.A(FE_OFN1809_acc_fir_data_in_0_));
   CLKINVX1TS FE_OFC1810_acc_fir_data_in_0_ (.Y(FE_OFN1810_acc_fir_data_in_0_), 
	.A(FE_OFN1809_acc_fir_data_in_0_));
   CLKINVX1TS FE_OFC1809_acc_fir_data_in_0_ (.Y(FE_OFN1809_acc_fir_data_in_0_), 
	.A(FE_OFN1808_acc_fir_data_in_0_));
   CLKBUFX2TS FE_OFC1808_acc_fir_data_in_0_ (.Y(FE_OFN1808_acc_fir_data_in_0_), 
	.A(acc_fir_data_in[0]));
   CLKBUFX2TS FE_OFC1807_acc_fir_data_in_1_ (.Y(FE_OFN1807_acc_fir_data_in_1_), 
	.A(FE_OFN1805_acc_fir_data_in_1_));
   CLKBUFX2TS FE_OFC1806_acc_fir_data_in_1_ (.Y(FE_OFN1806_acc_fir_data_in_1_), 
	.A(FE_OFN1805_acc_fir_data_in_1_));
   CLKBUFX2TS FE_OFC1805_acc_fir_data_in_1_ (.Y(FE_OFN1805_acc_fir_data_in_1_), 
	.A(FE_OFN1803_acc_fir_data_in_1_));
   CLKBUFX2TS FE_OFC1804_acc_fir_data_in_1_ (.Y(FE_OFN1804_acc_fir_data_in_1_), 
	.A(FE_OFN1803_acc_fir_data_in_1_));
   CLKBUFX2TS FE_OFC1803_acc_fir_data_in_1_ (.Y(FE_OFN1803_acc_fir_data_in_1_), 
	.A(FE_OFN1802_acc_fir_data_in_1_));
   CLKBUFX2TS FE_OFC1802_acc_fir_data_in_1_ (.Y(FE_OFN1802_acc_fir_data_in_1_), 
	.A(acc_fir_data_in[1]));
   CLKBUFX2TS FE_OFC1801_acc_fir_data_in_2_ (.Y(FE_OFN1801_acc_fir_data_in_2_), 
	.A(FE_OFN1800_acc_fir_data_in_2_));
   CLKINVX1TS FE_OFC1800_acc_fir_data_in_2_ (.Y(FE_OFN1800_acc_fir_data_in_2_), 
	.A(FE_OFN1798_acc_fir_data_in_2_));
   CLKINVX1TS FE_OFC1799_acc_fir_data_in_2_ (.Y(FE_OFN1799_acc_fir_data_in_2_), 
	.A(FE_OFN1798_acc_fir_data_in_2_));
   CLKINVX1TS FE_OFC1798_acc_fir_data_in_2_ (.Y(FE_OFN1798_acc_fir_data_in_2_), 
	.A(FE_OFN1797_acc_fir_data_in_2_));
   CLKBUFX2TS FE_OFC1797_acc_fir_data_in_2_ (.Y(FE_OFN1797_acc_fir_data_in_2_), 
	.A(FE_OFN1796_acc_fir_data_in_2_));
   CLKBUFX2TS FE_OFC1796_acc_fir_data_in_2_ (.Y(FE_OFN1796_acc_fir_data_in_2_), 
	.A(FE_OFN1795_acc_fir_data_in_2_));
   CLKBUFX2TS FE_OFC1795_acc_fir_data_in_2_ (.Y(FE_OFN1795_acc_fir_data_in_2_), 
	.A(acc_fir_data_in[2]));
   CLKBUFX2TS FE_OFC1794_acc_fir_data_in_3_ (.Y(FE_OFN1794_acc_fir_data_in_3_), 
	.A(FE_OFN1793_acc_fir_data_in_3_));
   CLKBUFX2TS FE_OFC1793_acc_fir_data_in_3_ (.Y(FE_OFN1793_acc_fir_data_in_3_), 
	.A(FE_OFN1791_acc_fir_data_in_3_));
   CLKBUFX2TS FE_OFC1792_acc_fir_data_in_3_ (.Y(FE_OFN1792_acc_fir_data_in_3_), 
	.A(FE_OFN1790_acc_fir_data_in_3_));
   CLKBUFX2TS FE_OFC1791_acc_fir_data_in_3_ (.Y(FE_OFN1791_acc_fir_data_in_3_), 
	.A(FE_OFN1790_acc_fir_data_in_3_));
   CLKBUFX2TS FE_OFC1790_acc_fir_data_in_3_ (.Y(FE_OFN1790_acc_fir_data_in_3_), 
	.A(acc_fir_data_in[3]));
   CLKBUFX2TS FE_OFC1789_acc_fir_data_in_4_ (.Y(FE_OFN1789_acc_fir_data_in_4_), 
	.A(FE_OFN1787_acc_fir_data_in_4_));
   CLKBUFX2TS FE_OFC1788_acc_fir_data_in_4_ (.Y(FE_OFN1788_acc_fir_data_in_4_), 
	.A(FE_OFN1786_acc_fir_data_in_4_));
   CLKBUFX2TS FE_OFC1787_acc_fir_data_in_4_ (.Y(FE_OFN1787_acc_fir_data_in_4_), 
	.A(FE_OFN1784_acc_fir_data_in_4_));
   CLKBUFX2TS FE_OFC1786_acc_fir_data_in_4_ (.Y(FE_OFN1786_acc_fir_data_in_4_), 
	.A(FE_OFN1785_acc_fir_data_in_4_));
   CLKINVX1TS FE_OFC1785_acc_fir_data_in_4_ (.Y(FE_OFN1785_acc_fir_data_in_4_), 
	.A(FE_OFN1783_acc_fir_data_in_4_));
   CLKINVX1TS FE_OFC1784_acc_fir_data_in_4_ (.Y(FE_OFN1784_acc_fir_data_in_4_), 
	.A(FE_OFN1783_acc_fir_data_in_4_));
   CLKINVX1TS FE_OFC1783_acc_fir_data_in_4_ (.Y(FE_OFN1783_acc_fir_data_in_4_), 
	.A(acc_fir_data_in[4]));
   CLKBUFX2TS FE_OFC1782_acc_fir_data_in_5_ (.Y(FE_OFN1782_acc_fir_data_in_5_), 
	.A(FE_OFN1781_acc_fir_data_in_5_));
   CLKBUFX2TS FE_OFC1781_acc_fir_data_in_5_ (.Y(FE_OFN1781_acc_fir_data_in_5_), 
	.A(FE_OFN1780_acc_fir_data_in_5_));
   CLKBUFX2TS FE_OFC1780_acc_fir_data_in_5_ (.Y(FE_OFN1780_acc_fir_data_in_5_), 
	.A(FE_OFN1778_acc_fir_data_in_5_));
   CLKBUFX2TS FE_OFC1779_acc_fir_data_in_5_ (.Y(FE_OFN1779_acc_fir_data_in_5_), 
	.A(FE_OFN1778_acc_fir_data_in_5_));
   CLKBUFX2TS FE_OFC1778_acc_fir_data_in_5_ (.Y(FE_OFN1778_acc_fir_data_in_5_), 
	.A(FE_OFN1777_acc_fir_data_in_5_));
   CLKBUFX2TS FE_OFC1777_acc_fir_data_in_5_ (.Y(FE_OFN1777_acc_fir_data_in_5_), 
	.A(acc_fir_data_in[5]));
   CLKBUFX2TS FE_OFC1776_acc_fir_data_in_6_ (.Y(FE_OFN1776_acc_fir_data_in_6_), 
	.A(FE_OFN1774_acc_fir_data_in_6_));
   CLKINVX1TS FE_OFC1775_acc_fir_data_in_6_ (.Y(FE_OFN1775_acc_fir_data_in_6_), 
	.A(FE_OFN1772_acc_fir_data_in_6_));
   CLKINVX1TS FE_OFC1774_acc_fir_data_in_6_ (.Y(FE_OFN1774_acc_fir_data_in_6_), 
	.A(FE_OFN1772_acc_fir_data_in_6_));
   CLKINVX1TS FE_OFC1773_acc_fir_data_in_6_ (.Y(FE_OFN1773_acc_fir_data_in_6_), 
	.A(FE_OFN1772_acc_fir_data_in_6_));
   CLKINVX1TS FE_OFC1772_acc_fir_data_in_6_ (.Y(FE_OFN1772_acc_fir_data_in_6_), 
	.A(FE_OFN1770_acc_fir_data_in_6_));
   CLKBUFX2TS FE_OFC1771_acc_fir_data_in_6_ (.Y(FE_OFN1771_acc_fir_data_in_6_), 
	.A(FE_OFN1770_acc_fir_data_in_6_));
   CLKBUFX2TS FE_OFC1770_acc_fir_data_in_6_ (.Y(FE_OFN1770_acc_fir_data_in_6_), 
	.A(FE_OFN1769_acc_fir_data_in_6_));
   CLKBUFX2TS FE_OFC1769_acc_fir_data_in_6_ (.Y(FE_OFN1769_acc_fir_data_in_6_), 
	.A(acc_fir_data_in[6]));
   CLKBUFX2TS FE_OFC1768_acc_fir_data_in_7_ (.Y(FE_OFN1768_acc_fir_data_in_7_), 
	.A(FE_OFN1765_acc_fir_data_in_7_));
   CLKBUFX2TS FE_OFC1767_acc_fir_data_in_7_ (.Y(FE_OFN1767_acc_fir_data_in_7_), 
	.A(FE_OFN1766_acc_fir_data_in_7_));
   CLKINVX1TS FE_OFC1766_acc_fir_data_in_7_ (.Y(FE_OFN1766_acc_fir_data_in_7_), 
	.A(FE_OFN1764_acc_fir_data_in_7_));
   CLKINVX1TS FE_OFC1765_acc_fir_data_in_7_ (.Y(FE_OFN1765_acc_fir_data_in_7_), 
	.A(FE_OFN1764_acc_fir_data_in_7_));
   INVX3TS FE_OFC1764_acc_fir_data_in_7_ (.Y(FE_OFN1764_acc_fir_data_in_7_), 
	.A(FE_OFN1763_acc_fir_data_in_7_));
   CLKBUFX2TS FE_OFC1763_acc_fir_data_in_7_ (.Y(FE_OFN1763_acc_fir_data_in_7_), 
	.A(FE_OFN1762_acc_fir_data_in_7_));
   CLKBUFX2TS FE_OFC1762_acc_fir_data_in_7_ (.Y(FE_OFN1762_acc_fir_data_in_7_), 
	.A(acc_fir_data_in[7]));
   CLKBUFX2TS FE_OFC1761_acc_fir_data_in_8_ (.Y(FE_OFN1761_acc_fir_data_in_8_), 
	.A(FE_OFN1759_acc_fir_data_in_8_));
   CLKBUFX2TS FE_OFC1760_acc_fir_data_in_8_ (.Y(FE_OFN1760_acc_fir_data_in_8_), 
	.A(FE_OFN1759_acc_fir_data_in_8_));
   CLKBUFX2TS FE_OFC1759_acc_fir_data_in_8_ (.Y(FE_OFN1759_acc_fir_data_in_8_), 
	.A(FE_OFN1758_acc_fir_data_in_8_));
   CLKBUFX2TS FE_OFC1758_acc_fir_data_in_8_ (.Y(FE_OFN1758_acc_fir_data_in_8_), 
	.A(FE_OFN1757_acc_fir_data_in_8_));
   CLKBUFX2TS FE_OFC1757_acc_fir_data_in_8_ (.Y(FE_OFN1757_acc_fir_data_in_8_), 
	.A(FE_OFN1756_acc_fir_data_in_8_));
   CLKBUFX2TS FE_OFC1756_acc_fir_data_in_8_ (.Y(FE_OFN1756_acc_fir_data_in_8_), 
	.A(acc_fir_data_in[8]));
   CLKBUFX2TS FE_OFC1755_acc_fir_data_in_9_ (.Y(FE_OFN1755_acc_fir_data_in_9_), 
	.A(FE_OFN1753_acc_fir_data_in_9_));
   CLKBUFX2TS FE_OFC1754_acc_fir_data_in_9_ (.Y(FE_OFN1754_acc_fir_data_in_9_), 
	.A(FE_OFN1752_acc_fir_data_in_9_));
   CLKBUFX2TS FE_OFC1753_acc_fir_data_in_9_ (.Y(FE_OFN1753_acc_fir_data_in_9_), 
	.A(FE_OFN1751_acc_fir_data_in_9_));
   CLKBUFX2TS FE_OFC1752_acc_fir_data_in_9_ (.Y(FE_OFN1752_acc_fir_data_in_9_), 
	.A(FE_OFN1751_acc_fir_data_in_9_));
   CLKBUFX2TS FE_OFC1751_acc_fir_data_in_9_ (.Y(FE_OFN1751_acc_fir_data_in_9_), 
	.A(acc_fir_data_in[9]));
   CLKBUFX2TS FE_OFC1750_acc_fir_data_in_10_ (.Y(FE_OFN1750_acc_fir_data_in_10_), 
	.A(FE_OFN1748_acc_fir_data_in_10_));
   CLKBUFX2TS FE_OFC1749_acc_fir_data_in_10_ (.Y(FE_OFN1749_acc_fir_data_in_10_), 
	.A(FE_OFN1747_acc_fir_data_in_10_));
   CLKBUFX2TS FE_OFC1748_acc_fir_data_in_10_ (.Y(FE_OFN1748_acc_fir_data_in_10_), 
	.A(FE_OFN1746_acc_fir_data_in_10_));
   CLKBUFX2TS FE_OFC1747_acc_fir_data_in_10_ (.Y(FE_OFN1747_acc_fir_data_in_10_), 
	.A(FE_OFN1746_acc_fir_data_in_10_));
   CLKBUFX2TS FE_OFC1746_acc_fir_data_in_10_ (.Y(FE_OFN1746_acc_fir_data_in_10_), 
	.A(acc_fir_data_in[10]));
   CLKBUFX2TS FE_OFC1745_acc_fir_data_in_11_ (.Y(FE_OFN1745_acc_fir_data_in_11_), 
	.A(FE_OFN1744_acc_fir_data_in_11_));
   CLKBUFX2TS FE_OFC1744_acc_fir_data_in_11_ (.Y(FE_OFN1744_acc_fir_data_in_11_), 
	.A(FE_OFN1743_acc_fir_data_in_11_));
   CLKBUFX2TS FE_OFC1743_acc_fir_data_in_11_ (.Y(FE_OFN1743_acc_fir_data_in_11_), 
	.A(FE_OFN1742_acc_fir_data_in_11_));
   CLKBUFX2TS FE_OFC1742_acc_fir_data_in_11_ (.Y(FE_OFN1742_acc_fir_data_in_11_), 
	.A(FE_OFN1741_acc_fir_data_in_11_));
   CLKBUFX2TS FE_OFC1741_acc_fir_data_in_11_ (.Y(FE_OFN1741_acc_fir_data_in_11_), 
	.A(acc_fir_data_in[11]));
   CLKBUFX2TS FE_OFC1740_acc_fir_data_in_12_ (.Y(FE_OFN1740_acc_fir_data_in_12_), 
	.A(FE_OFN1737_acc_fir_data_in_12_));
   CLKBUFX2TS FE_OFC1739_acc_fir_data_in_12_ (.Y(FE_OFN1739_acc_fir_data_in_12_), 
	.A(FE_OFN1738_acc_fir_data_in_12_));
   CLKBUFX2TS FE_OFC1738_acc_fir_data_in_12_ (.Y(FE_OFN1738_acc_fir_data_in_12_), 
	.A(FE_OFN1736_acc_fir_data_in_12_));
   CLKBUFX2TS FE_OFC1737_acc_fir_data_in_12_ (.Y(FE_OFN1737_acc_fir_data_in_12_), 
	.A(FE_OFN1736_acc_fir_data_in_12_));
   CLKBUFX2TS FE_OFC1736_acc_fir_data_in_12_ (.Y(FE_OFN1736_acc_fir_data_in_12_), 
	.A(acc_fir_data_in[12]));
   CLKBUFX2TS FE_OFC1735_acc_fir_data_in_13_ (.Y(FE_OFN1735_acc_fir_data_in_13_), 
	.A(FE_OFN1734_acc_fir_data_in_13_));
   CLKBUFX2TS FE_OFC1734_acc_fir_data_in_13_ (.Y(FE_OFN1734_acc_fir_data_in_13_), 
	.A(FE_OFN1733_acc_fir_data_in_13_));
   CLKBUFX2TS FE_OFC1733_acc_fir_data_in_13_ (.Y(FE_OFN1733_acc_fir_data_in_13_), 
	.A(FE_OFN1732_acc_fir_data_in_13_));
   CLKBUFX2TS FE_OFC1732_acc_fir_data_in_13_ (.Y(FE_OFN1732_acc_fir_data_in_13_), 
	.A(FE_OFN1731_acc_fir_data_in_13_));
   CLKBUFX2TS FE_OFC1731_acc_fir_data_in_13_ (.Y(FE_OFN1731_acc_fir_data_in_13_), 
	.A(acc_fir_data_in[13]));
   CLKBUFX2TS FE_OFC1730_acc_fir_data_in_14_ (.Y(FE_OFN1730_acc_fir_data_in_14_), 
	.A(FE_OFN1725_acc_fir_data_in_14_));
   CLKBUFX2TS FE_OFC1729_acc_fir_data_in_14_ (.Y(FE_OFN1729_acc_fir_data_in_14_), 
	.A(FE_OFN1727_acc_fir_data_in_14_));
   CLKINVX1TS FE_OFC1728_acc_fir_data_in_14_ (.Y(FE_OFN1728_acc_fir_data_in_14_), 
	.A(FE_OFN1726_acc_fir_data_in_14_));
   CLKINVX1TS FE_OFC1727_acc_fir_data_in_14_ (.Y(FE_OFN1727_acc_fir_data_in_14_), 
	.A(FE_OFN1726_acc_fir_data_in_14_));
   CLKINVX1TS FE_OFC1726_acc_fir_data_in_14_ (.Y(FE_OFN1726_acc_fir_data_in_14_), 
	.A(FE_OFN1724_acc_fir_data_in_14_));
   CLKBUFX2TS FE_OFC1725_acc_fir_data_in_14_ (.Y(FE_OFN1725_acc_fir_data_in_14_), 
	.A(FE_OFN1724_acc_fir_data_in_14_));
   CLKBUFX2TS FE_OFC1724_acc_fir_data_in_14_ (.Y(FE_OFN1724_acc_fir_data_in_14_), 
	.A(acc_fir_data_in[14]));
   CLKBUFX2TS FE_OFC1723_acc_fir_data_in_15_ (.Y(FE_OFN1723_acc_fir_data_in_15_), 
	.A(FE_OFN1720_acc_fir_data_in_15_));
   CLKBUFX2TS FE_OFC1722_acc_fir_data_in_15_ (.Y(FE_OFN1722_acc_fir_data_in_15_), 
	.A(FE_OFN1721_acc_fir_data_in_15_));
   CLKBUFX2TS FE_OFC1721_acc_fir_data_in_15_ (.Y(FE_OFN1721_acc_fir_data_in_15_), 
	.A(FE_OFN1719_acc_fir_data_in_15_));
   CLKBUFX2TS FE_OFC1720_acc_fir_data_in_15_ (.Y(FE_OFN1720_acc_fir_data_in_15_), 
	.A(FE_OFN1719_acc_fir_data_in_15_));
   CLKBUFX2TS FE_OFC1719_acc_fir_data_in_15_ (.Y(FE_OFN1719_acc_fir_data_in_15_), 
	.A(acc_fir_data_in[15]));
   CLKBUFX2TS FE_OFC1718_acc_fir_data_in_16_ (.Y(FE_OFN1718_acc_fir_data_in_16_), 
	.A(FE_OFN1717_acc_fir_data_in_16_));
   CLKBUFX2TS FE_OFC1717_acc_fir_data_in_16_ (.Y(FE_OFN1717_acc_fir_data_in_16_), 
	.A(FE_OFN1715_acc_fir_data_in_16_));
   CLKINVX1TS FE_OFC1716_acc_fir_data_in_16_ (.Y(FE_OFN1716_acc_fir_data_in_16_), 
	.A(FE_OFN1714_acc_fir_data_in_16_));
   CLKINVX1TS FE_OFC1715_acc_fir_data_in_16_ (.Y(FE_OFN1715_acc_fir_data_in_16_), 
	.A(FE_OFN1714_acc_fir_data_in_16_));
   CLKINVX1TS FE_OFC1714_acc_fir_data_in_16_ (.Y(FE_OFN1714_acc_fir_data_in_16_), 
	.A(FE_OFN1713_acc_fir_data_in_16_));
   CLKBUFX2TS FE_OFC1713_acc_fir_data_in_16_ (.Y(FE_OFN1713_acc_fir_data_in_16_), 
	.A(FE_OFN1712_acc_fir_data_in_16_));
   CLKBUFX2TS FE_OFC1712_acc_fir_data_in_16_ (.Y(FE_OFN1712_acc_fir_data_in_16_), 
	.A(acc_fir_data_in[16]));
   CLKBUFX2TS FE_OFC1711_acc_fir_data_in_17_ (.Y(FE_OFN1711_acc_fir_data_in_17_), 
	.A(FE_OFN1708_acc_fir_data_in_17_));
   CLKBUFX2TS FE_OFC1710_acc_fir_data_in_17_ (.Y(FE_OFN1710_acc_fir_data_in_17_), 
	.A(FE_OFN1709_acc_fir_data_in_17_));
   CLKBUFX2TS FE_OFC1709_acc_fir_data_in_17_ (.Y(FE_OFN1709_acc_fir_data_in_17_), 
	.A(FE_OFN1707_acc_fir_data_in_17_));
   CLKBUFX2TS FE_OFC1708_acc_fir_data_in_17_ (.Y(FE_OFN1708_acc_fir_data_in_17_), 
	.A(FE_OFN1707_acc_fir_data_in_17_));
   CLKBUFX2TS FE_OFC1707_acc_fir_data_in_17_ (.Y(FE_OFN1707_acc_fir_data_in_17_), 
	.A(acc_fir_data_in[17]));
   CLKBUFX2TS FE_OFC1706_acc_fir_data_in_18_ (.Y(FE_OFN1706_acc_fir_data_in_18_), 
	.A(FE_OFN1705_acc_fir_data_in_18_));
   CLKBUFX2TS FE_OFC1705_acc_fir_data_in_18_ (.Y(FE_OFN1705_acc_fir_data_in_18_), 
	.A(FE_OFN1704_acc_fir_data_in_18_));
   CLKBUFX2TS FE_OFC1704_acc_fir_data_in_18_ (.Y(FE_OFN1704_acc_fir_data_in_18_), 
	.A(FE_OFN1703_acc_fir_data_in_18_));
   CLKBUFX2TS FE_OFC1703_acc_fir_data_in_18_ (.Y(FE_OFN1703_acc_fir_data_in_18_), 
	.A(FE_OFN1702_acc_fir_data_in_18_));
   CLKBUFX2TS FE_OFC1702_acc_fir_data_in_18_ (.Y(FE_OFN1702_acc_fir_data_in_18_), 
	.A(acc_fir_data_in[18]));
   CLKBUFX2TS FE_OFC1701_acc_fir_data_in_19_ (.Y(FE_OFN1701_acc_fir_data_in_19_), 
	.A(FE_OFN1699_acc_fir_data_in_19_));
   CLKBUFX2TS FE_OFC1700_acc_fir_data_in_19_ (.Y(FE_OFN1700_acc_fir_data_in_19_), 
	.A(FE_OFN1699_acc_fir_data_in_19_));
   CLKBUFX2TS FE_OFC1699_acc_fir_data_in_19_ (.Y(FE_OFN1699_acc_fir_data_in_19_), 
	.A(FE_OFN1698_acc_fir_data_in_19_));
   CLKINVX1TS FE_OFC1698_acc_fir_data_in_19_ (.Y(FE_OFN1698_acc_fir_data_in_19_), 
	.A(FE_OFN1696_acc_fir_data_in_19_));
   CLKINVX1TS FE_OFC1697_acc_fir_data_in_19_ (.Y(FE_OFN1697_acc_fir_data_in_19_), 
	.A(FE_OFN1696_acc_fir_data_in_19_));
   CLKINVX1TS FE_OFC1696_acc_fir_data_in_19_ (.Y(FE_OFN1696_acc_fir_data_in_19_), 
	.A(FE_OFN1695_acc_fir_data_in_19_));
   CLKBUFX2TS FE_OFC1695_acc_fir_data_in_19_ (.Y(FE_OFN1695_acc_fir_data_in_19_), 
	.A(acc_fir_data_in[19]));
   CLKBUFX2TS FE_OFC1694_acc_fir_data_in_20_ (.Y(FE_OFN1694_acc_fir_data_in_20_), 
	.A(FE_OFN1692_acc_fir_data_in_20_));
   CLKBUFX2TS FE_OFC1693_acc_fir_data_in_20_ (.Y(FE_OFN1693_acc_fir_data_in_20_), 
	.A(FE_OFN1691_acc_fir_data_in_20_));
   CLKBUFX2TS FE_OFC1692_acc_fir_data_in_20_ (.Y(FE_OFN1692_acc_fir_data_in_20_), 
	.A(FE_OFN1691_acc_fir_data_in_20_));
   CLKBUFX2TS FE_OFC1691_acc_fir_data_in_20_ (.Y(FE_OFN1691_acc_fir_data_in_20_), 
	.A(FE_OFN1690_acc_fir_data_in_20_));
   CLKBUFX2TS FE_OFC1690_acc_fir_data_in_20_ (.Y(FE_OFN1690_acc_fir_data_in_20_), 
	.A(acc_fir_data_in[20]));
   CLKBUFX2TS FE_OFC1689_acc_fir_data_in_21_ (.Y(FE_OFN1689_acc_fir_data_in_21_), 
	.A(FE_OFN1687_acc_fir_data_in_21_));
   CLKINVX1TS FE_OFC1688_acc_fir_data_in_21_ (.Y(FE_OFN1688_acc_fir_data_in_21_), 
	.A(FE_OFN1686_acc_fir_data_in_21_));
   CLKINVX1TS FE_OFC1687_acc_fir_data_in_21_ (.Y(FE_OFN1687_acc_fir_data_in_21_), 
	.A(FE_OFN1686_acc_fir_data_in_21_));
   CLKINVX1TS FE_OFC1686_acc_fir_data_in_21_ (.Y(FE_OFN1686_acc_fir_data_in_21_), 
	.A(FE_OFN1685_acc_fir_data_in_21_));
   CLKBUFX2TS FE_OFC1685_acc_fir_data_in_21_ (.Y(FE_OFN1685_acc_fir_data_in_21_), 
	.A(FE_OFN1684_acc_fir_data_in_21_));
   CLKBUFX2TS FE_OFC1684_acc_fir_data_in_21_ (.Y(FE_OFN1684_acc_fir_data_in_21_), 
	.A(FE_OFN1683_acc_fir_data_in_21_));
   CLKBUFX2TS FE_OFC1683_acc_fir_data_in_21_ (.Y(FE_OFN1683_acc_fir_data_in_21_), 
	.A(acc_fir_data_in[21]));
   CLKBUFX2TS FE_OFC1682_acc_fir_data_in_22_ (.Y(FE_OFN1682_acc_fir_data_in_22_), 
	.A(FE_OFN1681_acc_fir_data_in_22_));
   CLKBUFX2TS FE_OFC1681_acc_fir_data_in_22_ (.Y(FE_OFN1681_acc_fir_data_in_22_), 
	.A(FE_OFN1680_acc_fir_data_in_22_));
   CLKBUFX2TS FE_OFC1680_acc_fir_data_in_22_ (.Y(FE_OFN1680_acc_fir_data_in_22_), 
	.A(FE_OFN1678_acc_fir_data_in_22_));
   CLKBUFX2TS FE_OFC1679_acc_fir_data_in_22_ (.Y(FE_OFN1679_acc_fir_data_in_22_), 
	.A(FE_OFN1678_acc_fir_data_in_22_));
   CLKBUFX2TS FE_OFC1678_acc_fir_data_in_22_ (.Y(FE_OFN1678_acc_fir_data_in_22_), 
	.A(acc_fir_data_in[22]));
   CLKBUFX2TS FE_OFC1677_acc_fir_data_in_23_ (.Y(FE_OFN1677_acc_fir_data_in_23_), 
	.A(FE_OFN1675_acc_fir_data_in_23_));
   CLKINVX1TS FE_OFC1676_acc_fir_data_in_23_ (.Y(FE_OFN1676_acc_fir_data_in_23_), 
	.A(FE_OFN1674_acc_fir_data_in_23_));
   CLKINVX1TS FE_OFC1675_acc_fir_data_in_23_ (.Y(FE_OFN1675_acc_fir_data_in_23_), 
	.A(FE_OFN1674_acc_fir_data_in_23_));
   CLKINVX1TS FE_OFC1674_acc_fir_data_in_23_ (.Y(FE_OFN1674_acc_fir_data_in_23_), 
	.A(FE_OFN1672_acc_fir_data_in_23_));
   CLKBUFX2TS FE_OFC1673_acc_fir_data_in_23_ (.Y(FE_OFN1673_acc_fir_data_in_23_), 
	.A(FE_OFN1672_acc_fir_data_in_23_));
   CLKBUFX2TS FE_OFC1672_acc_fir_data_in_23_ (.Y(FE_OFN1672_acc_fir_data_in_23_), 
	.A(FE_OFN1671_acc_fir_data_in_23_));
   CLKBUFX2TS FE_OFC1671_acc_fir_data_in_23_ (.Y(FE_OFN1671_acc_fir_data_in_23_), 
	.A(acc_fir_data_in[23]));
   CLKBUFX2TS FE_OFC1670_acc_fir_data_in_24_ (.Y(FE_OFN1670_acc_fir_data_in_24_), 
	.A(FE_OFN1669_acc_fir_data_in_24_));
   CLKBUFX2TS FE_OFC1669_acc_fir_data_in_24_ (.Y(FE_OFN1669_acc_fir_data_in_24_), 
	.A(FE_OFN1667_acc_fir_data_in_24_));
   CLKBUFX2TS FE_OFC1668_acc_fir_data_in_24_ (.Y(FE_OFN1668_acc_fir_data_in_24_), 
	.A(FE_OFN1667_acc_fir_data_in_24_));
   CLKBUFX2TS FE_OFC1667_acc_fir_data_in_24_ (.Y(FE_OFN1667_acc_fir_data_in_24_), 
	.A(FE_OFN1666_acc_fir_data_in_24_));
   CLKBUFX2TS FE_OFC1666_acc_fir_data_in_24_ (.Y(FE_OFN1666_acc_fir_data_in_24_), 
	.A(acc_fir_data_in[24]));
   CLKBUFX2TS FE_OFC1665_acc_fir_data_in_25_ (.Y(FE_OFN1665_acc_fir_data_in_25_), 
	.A(FE_OFN1664_acc_fir_data_in_25_));
   CLKBUFX2TS FE_OFC1664_acc_fir_data_in_25_ (.Y(FE_OFN1664_acc_fir_data_in_25_), 
	.A(FE_OFN1663_acc_fir_data_in_25_));
   CLKBUFX2TS FE_OFC1663_acc_fir_data_in_25_ (.Y(FE_OFN1663_acc_fir_data_in_25_), 
	.A(FE_OFN1662_acc_fir_data_in_25_));
   CLKBUFX2TS FE_OFC1662_acc_fir_data_in_25_ (.Y(FE_OFN1662_acc_fir_data_in_25_), 
	.A(FE_OFN1661_acc_fir_data_in_25_));
   CLKBUFX2TS FE_OFC1661_acc_fir_data_in_25_ (.Y(FE_OFN1661_acc_fir_data_in_25_), 
	.A(acc_fir_data_in[25]));
   CLKBUFX2TS FE_OFC1660_acc_fir_data_in_26_ (.Y(FE_OFN1660_acc_fir_data_in_26_), 
	.A(FE_OFN1659_acc_fir_data_in_26_));
   CLKBUFX2TS FE_OFC1659_acc_fir_data_in_26_ (.Y(FE_OFN1659_acc_fir_data_in_26_), 
	.A(FE_OFN1818_acc_fir_data_in_26_));
   CLKBUFX2TS FE_OFC1658_acc_fir_data_in_26_ (.Y(FE_OFN1658_acc_fir_data_in_26_), 
	.A(FE_OFN1657_acc_fir_data_in_26_));
   CLKBUFX2TS FE_OFC1657_acc_fir_data_in_26_ (.Y(FE_OFN1657_acc_fir_data_in_26_), 
	.A(FE_OFN1818_acc_fir_data_in_26_));
   CLKBUFX2TS FE_OFC1656_acc_fir_data_in_26_ (.Y(FE_OFN1656_acc_fir_data_in_26_), 
	.A(acc_fir_data_in[26]));
   CLKBUFX2TS FE_OFC1655_acc_fir_data_in_27_ (.Y(FE_OFN1655_acc_fir_data_in_27_), 
	.A(FE_OFN1653_acc_fir_data_in_27_));
   CLKBUFX2TS FE_OFC1654_acc_fir_data_in_27_ (.Y(FE_OFN1654_acc_fir_data_in_27_), 
	.A(FE_OFN1652_acc_fir_data_in_27_));
   CLKBUFX2TS FE_OFC1653_acc_fir_data_in_27_ (.Y(FE_OFN1653_acc_fir_data_in_27_), 
	.A(FE_OFN1651_acc_fir_data_in_27_));
   CLKBUFX2TS FE_OFC1652_acc_fir_data_in_27_ (.Y(FE_OFN1652_acc_fir_data_in_27_), 
	.A(FE_OFN1651_acc_fir_data_in_27_));
   CLKBUFX2TS FE_OFC1651_acc_fir_data_in_27_ (.Y(FE_OFN1651_acc_fir_data_in_27_), 
	.A(acc_fir_data_in[27]));
   CLKBUFX2TS FE_OFC1650_acc_fir_data_in_28_ (.Y(FE_OFN1650_acc_fir_data_in_28_), 
	.A(FE_OFN1648_acc_fir_data_in_28_));
   CLKBUFX2TS FE_OFC1649_acc_fir_data_in_28_ (.Y(FE_OFN1649_acc_fir_data_in_28_), 
	.A(FE_OFN1647_acc_fir_data_in_28_));
   CLKBUFX2TS FE_OFC1648_acc_fir_data_in_28_ (.Y(FE_OFN1648_acc_fir_data_in_28_), 
	.A(FE_OFN1646_acc_fir_data_in_28_));
   CLKBUFX2TS FE_OFC1647_acc_fir_data_in_28_ (.Y(FE_OFN1647_acc_fir_data_in_28_), 
	.A(FE_OFN1646_acc_fir_data_in_28_));
   CLKBUFX2TS FE_OFC1646_acc_fir_data_in_28_ (.Y(FE_OFN1646_acc_fir_data_in_28_), 
	.A(acc_fir_data_in[28]));
   CLKBUFX2TS FE_OFC1645_acc_fir_data_in_29_ (.Y(FE_OFN1645_acc_fir_data_in_29_), 
	.A(FE_OFN1643_acc_fir_data_in_29_));
   CLKBUFX2TS FE_OFC1644_acc_fir_data_in_29_ (.Y(FE_OFN1644_acc_fir_data_in_29_), 
	.A(FE_OFN1643_acc_fir_data_in_29_));
   CLKBUFX2TS FE_OFC1643_acc_fir_data_in_29_ (.Y(FE_OFN1643_acc_fir_data_in_29_), 
	.A(FE_OFN1641_acc_fir_data_in_29_));
   CLKINVX1TS FE_OFC1642_acc_fir_data_in_29_ (.Y(FE_OFN1642_acc_fir_data_in_29_), 
	.A(FE_OFN1639_acc_fir_data_in_29_));
   CLKINVX1TS FE_OFC1641_acc_fir_data_in_29_ (.Y(FE_OFN1641_acc_fir_data_in_29_), 
	.A(FE_OFN1639_acc_fir_data_in_29_));
   CLKINVX1TS FE_OFC1640_acc_fir_data_in_29_ (.Y(FE_OFN1640_acc_fir_data_in_29_), 
	.A(FE_OFN1639_acc_fir_data_in_29_));
   CLKINVX1TS FE_OFC1639_acc_fir_data_in_29_ (.Y(FE_OFN1639_acc_fir_data_in_29_), 
	.A(FE_OFN1638_acc_fir_data_in_29_));
   CLKBUFX2TS FE_OFC1638_acc_fir_data_in_29_ (.Y(FE_OFN1638_acc_fir_data_in_29_), 
	.A(acc_fir_data_in[29]));
   CLKBUFX2TS FE_OFC1637_acc_fir_data_in_30_ (.Y(FE_OFN1637_acc_fir_data_in_30_), 
	.A(FE_OFN1635_acc_fir_data_in_30_));
   CLKBUFX2TS FE_OFC1636_acc_fir_data_in_30_ (.Y(FE_OFN1636_acc_fir_data_in_30_), 
	.A(FE_OFN1634_acc_fir_data_in_30_));
   CLKBUFX2TS FE_OFC1635_acc_fir_data_in_30_ (.Y(FE_OFN1635_acc_fir_data_in_30_), 
	.A(FE_OFN1633_acc_fir_data_in_30_));
   CLKBUFX2TS FE_OFC1634_acc_fir_data_in_30_ (.Y(FE_OFN1634_acc_fir_data_in_30_), 
	.A(FE_OFN1633_acc_fir_data_in_30_));
   CLKBUFX2TS FE_OFC1633_acc_fir_data_in_30_ (.Y(FE_OFN1633_acc_fir_data_in_30_), 
	.A(acc_fir_data_in[30]));
   CLKBUFX2TS FE_OFC1632_acc_fir_data_in_31_ (.Y(FE_OFN1632_acc_fir_data_in_31_), 
	.A(FE_OFN1630_acc_fir_data_in_31_));
   CLKBUFX2TS FE_OFC1631_acc_fir_data_in_31_ (.Y(FE_OFN1631_acc_fir_data_in_31_), 
	.A(FE_OFN1630_acc_fir_data_in_31_));
   CLKBUFX2TS FE_OFC1630_acc_fir_data_in_31_ (.Y(FE_OFN1630_acc_fir_data_in_31_), 
	.A(FE_OFN1629_acc_fir_data_in_31_));
   CLKBUFX2TS FE_OFC1629_acc_fir_data_in_31_ (.Y(FE_OFN1629_acc_fir_data_in_31_), 
	.A(FE_OFN1628_acc_fir_data_in_31_));
   CLKBUFX2TS FE_OFC1628_acc_fir_data_in_31_ (.Y(FE_OFN1628_acc_fir_data_in_31_), 
	.A(acc_fir_data_in[31]));
   CLKBUFX2TS FE_OFC1627_acc_fft_data_in_0_ (.Y(FE_OFN1627_acc_fft_data_in_0_), 
	.A(FE_OFN1626_acc_fft_data_in_0_));
   CLKBUFX2TS FE_OFC1626_acc_fft_data_in_0_ (.Y(FE_OFN1626_acc_fft_data_in_0_), 
	.A(FE_OFN1625_acc_fft_data_in_0_));
   CLKBUFX2TS FE_OFC1625_acc_fft_data_in_0_ (.Y(FE_OFN1625_acc_fft_data_in_0_), 
	.A(FE_OFN1624_acc_fft_data_in_0_));
   CLKBUFX2TS FE_OFC1624_acc_fft_data_in_0_ (.Y(FE_OFN1624_acc_fft_data_in_0_), 
	.A(FE_OFN1623_acc_fft_data_in_0_));
   CLKBUFX2TS FE_OFC1623_acc_fft_data_in_0_ (.Y(FE_OFN1623_acc_fft_data_in_0_), 
	.A(FE_OFN1622_acc_fft_data_in_0_));
   CLKBUFX2TS FE_OFC1622_acc_fft_data_in_0_ (.Y(FE_OFN1622_acc_fft_data_in_0_), 
	.A(acc_fft_data_in[0]));
   CLKINVX1TS FE_OFC1621_acc_fft_data_in_1_ (.Y(FE_OFN1621_acc_fft_data_in_1_), 
	.A(FE_OFN1619_acc_fft_data_in_1_));
   CLKINVX1TS FE_OFC1620_acc_fft_data_in_1_ (.Y(FE_OFN1620_acc_fft_data_in_1_), 
	.A(FE_OFN1619_acc_fft_data_in_1_));
   CLKINVX1TS FE_OFC1619_acc_fft_data_in_1_ (.Y(FE_OFN1619_acc_fft_data_in_1_), 
	.A(FE_OFN1618_acc_fft_data_in_1_));
   CLKBUFX2TS FE_OFC1618_acc_fft_data_in_1_ (.Y(FE_OFN1618_acc_fft_data_in_1_), 
	.A(FE_OFN1617_acc_fft_data_in_1_));
   CLKBUFX2TS FE_OFC1617_acc_fft_data_in_1_ (.Y(FE_OFN1617_acc_fft_data_in_1_), 
	.A(FE_OFN1616_acc_fft_data_in_1_));
   CLKBUFX2TS FE_OFC1616_acc_fft_data_in_1_ (.Y(FE_OFN1616_acc_fft_data_in_1_), 
	.A(FE_OFN1615_acc_fft_data_in_1_));
   CLKBUFX2TS FE_OFC1615_acc_fft_data_in_1_ (.Y(FE_OFN1615_acc_fft_data_in_1_), 
	.A(acc_fft_data_in[1]));
   CLKBUFX2TS FE_OFC1614_acc_fft_data_in_2_ (.Y(FE_OFN1614_acc_fft_data_in_2_), 
	.A(FE_OFN1612_acc_fft_data_in_2_));
   CLKINVX1TS FE_OFC1613_acc_fft_data_in_2_ (.Y(FE_OFN1613_acc_fft_data_in_2_), 
	.A(FE_OFN1611_acc_fft_data_in_2_));
   CLKINVX1TS FE_OFC1612_acc_fft_data_in_2_ (.Y(FE_OFN1612_acc_fft_data_in_2_), 
	.A(FE_OFN1611_acc_fft_data_in_2_));
   CLKINVX1TS FE_OFC1611_acc_fft_data_in_2_ (.Y(FE_OFN1611_acc_fft_data_in_2_), 
	.A(FE_OFN1610_acc_fft_data_in_2_));
   CLKBUFX2TS FE_OFC1610_acc_fft_data_in_2_ (.Y(FE_OFN1610_acc_fft_data_in_2_), 
	.A(FE_OFN1609_acc_fft_data_in_2_));
   CLKBUFX2TS FE_OFC1609_acc_fft_data_in_2_ (.Y(FE_OFN1609_acc_fft_data_in_2_), 
	.A(FE_OFN1608_acc_fft_data_in_2_));
   CLKBUFX2TS FE_OFC1608_acc_fft_data_in_2_ (.Y(FE_OFN1608_acc_fft_data_in_2_), 
	.A(acc_fft_data_in[2]));
   CLKBUFX2TS FE_OFC1607_acc_fft_data_in_3_ (.Y(FE_OFN1607_acc_fft_data_in_3_), 
	.A(FE_OFN1605_acc_fft_data_in_3_));
   CLKBUFX2TS FE_OFC1606_acc_fft_data_in_3_ (.Y(FE_OFN1606_acc_fft_data_in_3_), 
	.A(FE_OFN1605_acc_fft_data_in_3_));
   CLKBUFX2TS FE_OFC1605_acc_fft_data_in_3_ (.Y(FE_OFN1605_acc_fft_data_in_3_), 
	.A(FE_OFN1604_acc_fft_data_in_3_));
   CLKBUFX2TS FE_OFC1604_acc_fft_data_in_3_ (.Y(FE_OFN1604_acc_fft_data_in_3_), 
	.A(FE_OFN1603_acc_fft_data_in_3_));
   CLKBUFX2TS FE_OFC1603_acc_fft_data_in_3_ (.Y(FE_OFN1603_acc_fft_data_in_3_), 
	.A(acc_fft_data_in[3]));
   CLKBUFX2TS FE_OFC1602_acc_fft_data_in_4_ (.Y(FE_OFN1602_acc_fft_data_in_4_), 
	.A(FE_OFN1601_acc_fft_data_in_4_));
   CLKBUFX2TS FE_OFC1601_acc_fft_data_in_4_ (.Y(FE_OFN1601_acc_fft_data_in_4_), 
	.A(FE_OFN1600_acc_fft_data_in_4_));
   CLKBUFX2TS FE_OFC1600_acc_fft_data_in_4_ (.Y(FE_OFN1600_acc_fft_data_in_4_), 
	.A(FE_OFN1597_acc_fft_data_in_4_));
   CLKBUFX2TS FE_OFC1599_acc_fft_data_in_4_ (.Y(FE_OFN1599_acc_fft_data_in_4_), 
	.A(FE_OFN1598_acc_fft_data_in_4_));
   CLKINVX1TS FE_OFC1598_acc_fft_data_in_4_ (.Y(FE_OFN1598_acc_fft_data_in_4_), 
	.A(FE_OFN1596_acc_fft_data_in_4_));
   CLKINVX1TS FE_OFC1597_acc_fft_data_in_4_ (.Y(FE_OFN1597_acc_fft_data_in_4_), 
	.A(FE_OFN1596_acc_fft_data_in_4_));
   CLKINVX2TS FE_OFC1596_acc_fft_data_in_4_ (.Y(FE_OFN1596_acc_fft_data_in_4_), 
	.A(acc_fft_data_in[4]));
   CLKBUFX2TS FE_OFC1595_acc_fft_data_in_5_ (.Y(FE_OFN1595_acc_fft_data_in_5_), 
	.A(FE_OFN1593_acc_fft_data_in_5_));
   CLKBUFX2TS FE_OFC1594_acc_fft_data_in_5_ (.Y(FE_OFN1594_acc_fft_data_in_5_), 
	.A(FE_OFN1592_acc_fft_data_in_5_));
   CLKBUFX2TS FE_OFC1593_acc_fft_data_in_5_ (.Y(FE_OFN1593_acc_fft_data_in_5_), 
	.A(FE_OFN1592_acc_fft_data_in_5_));
   CLKBUFX2TS FE_OFC1592_acc_fft_data_in_5_ (.Y(FE_OFN1592_acc_fft_data_in_5_), 
	.A(FE_OFN1591_acc_fft_data_in_5_));
   CLKBUFX2TS FE_OFC1591_acc_fft_data_in_5_ (.Y(FE_OFN1591_acc_fft_data_in_5_), 
	.A(acc_fft_data_in[5]));
   CLKBUFX2TS FE_OFC1590_acc_fft_data_in_6_ (.Y(FE_OFN1590_acc_fft_data_in_6_), 
	.A(FE_OFN1588_acc_fft_data_in_6_));
   CLKBUFX2TS FE_OFC1589_acc_fft_data_in_6_ (.Y(FE_OFN1589_acc_fft_data_in_6_), 
	.A(FE_OFN1588_acc_fft_data_in_6_));
   CLKBUFX2TS FE_OFC1588_acc_fft_data_in_6_ (.Y(FE_OFN1588_acc_fft_data_in_6_), 
	.A(FE_OFN1587_acc_fft_data_in_6_));
   CLKBUFX2TS FE_OFC1587_acc_fft_data_in_6_ (.Y(FE_OFN1587_acc_fft_data_in_6_), 
	.A(FE_OFN1586_acc_fft_data_in_6_));
   CLKBUFX2TS FE_OFC1586_acc_fft_data_in_6_ (.Y(FE_OFN1586_acc_fft_data_in_6_), 
	.A(FE_OFN1585_acc_fft_data_in_6_));
   CLKBUFX2TS FE_OFC1585_acc_fft_data_in_6_ (.Y(FE_OFN1585_acc_fft_data_in_6_), 
	.A(acc_fft_data_in[6]));
   CLKBUFX2TS FE_OFC1584_acc_fft_data_in_7_ (.Y(FE_OFN1584_acc_fft_data_in_7_), 
	.A(FE_OFN1583_acc_fft_data_in_7_));
   CLKBUFX2TS FE_OFC1583_acc_fft_data_in_7_ (.Y(FE_OFN1583_acc_fft_data_in_7_), 
	.A(FE_OFN1582_acc_fft_data_in_7_));
   CLKBUFX2TS FE_OFC1582_acc_fft_data_in_7_ (.Y(FE_OFN1582_acc_fft_data_in_7_), 
	.A(FE_OFN1580_acc_fft_data_in_7_));
   CLKBUFX2TS FE_OFC1581_acc_fft_data_in_7_ (.Y(FE_OFN1581_acc_fft_data_in_7_), 
	.A(FE_OFN1580_acc_fft_data_in_7_));
   CLKBUFX2TS FE_OFC1580_acc_fft_data_in_7_ (.Y(FE_OFN1580_acc_fft_data_in_7_), 
	.A(acc_fft_data_in[7]));
   CLKBUFX2TS FE_OFC1579_acc_fft_data_in_8_ (.Y(FE_OFN1579_acc_fft_data_in_8_), 
	.A(FE_OFN1578_acc_fft_data_in_8_));
   CLKBUFX2TS FE_OFC1578_acc_fft_data_in_8_ (.Y(FE_OFN1578_acc_fft_data_in_8_), 
	.A(FE_OFN1577_acc_fft_data_in_8_));
   CLKBUFX2TS FE_OFC1577_acc_fft_data_in_8_ (.Y(FE_OFN1577_acc_fft_data_in_8_), 
	.A(FE_OFN1576_acc_fft_data_in_8_));
   CLKBUFX2TS FE_OFC1576_acc_fft_data_in_8_ (.Y(FE_OFN1576_acc_fft_data_in_8_), 
	.A(FE_OFN1575_acc_fft_data_in_8_));
   CLKBUFX2TS FE_OFC1575_acc_fft_data_in_8_ (.Y(FE_OFN1575_acc_fft_data_in_8_), 
	.A(FE_OFN1574_acc_fft_data_in_8_));
   CLKBUFX2TS FE_OFC1574_acc_fft_data_in_8_ (.Y(FE_OFN1574_acc_fft_data_in_8_), 
	.A(acc_fft_data_in[8]));
   CLKBUFX2TS FE_OFC1573_acc_fft_data_in_9_ (.Y(FE_OFN1573_acc_fft_data_in_9_), 
	.A(FE_OFN1571_acc_fft_data_in_9_));
   CLKBUFX2TS FE_OFC1572_acc_fft_data_in_9_ (.Y(FE_OFN1572_acc_fft_data_in_9_), 
	.A(FE_OFN1570_acc_fft_data_in_9_));
   CLKBUFX2TS FE_OFC1571_acc_fft_data_in_9_ (.Y(FE_OFN1571_acc_fft_data_in_9_), 
	.A(FE_OFN1569_acc_fft_data_in_9_));
   CLKBUFX2TS FE_OFC1570_acc_fft_data_in_9_ (.Y(FE_OFN1570_acc_fft_data_in_9_), 
	.A(FE_OFN1569_acc_fft_data_in_9_));
   CLKBUFX2TS FE_OFC1569_acc_fft_data_in_9_ (.Y(FE_OFN1569_acc_fft_data_in_9_), 
	.A(acc_fft_data_in[9]));
   CLKBUFX2TS FE_OFC1568_acc_fft_data_in_10_ (.Y(FE_OFN1568_acc_fft_data_in_10_), 
	.A(FE_OFN1565_acc_fft_data_in_10_));
   CLKBUFX2TS FE_OFC1567_acc_fft_data_in_10_ (.Y(FE_OFN1567_acc_fft_data_in_10_), 
	.A(FE_OFN1566_acc_fft_data_in_10_));
   CLKBUFX2TS FE_OFC1566_acc_fft_data_in_10_ (.Y(FE_OFN1566_acc_fft_data_in_10_), 
	.A(FE_OFN1564_acc_fft_data_in_10_));
   CLKBUFX2TS FE_OFC1565_acc_fft_data_in_10_ (.Y(FE_OFN1565_acc_fft_data_in_10_), 
	.A(FE_OFN1564_acc_fft_data_in_10_));
   CLKBUFX2TS FE_OFC1564_acc_fft_data_in_10_ (.Y(FE_OFN1564_acc_fft_data_in_10_), 
	.A(acc_fft_data_in[10]));
   CLKBUFX2TS FE_OFC1563_acc_fft_data_in_11_ (.Y(FE_OFN1563_acc_fft_data_in_11_), 
	.A(FE_OFN1562_acc_fft_data_in_11_));
   CLKBUFX2TS FE_OFC1562_acc_fft_data_in_11_ (.Y(FE_OFN1562_acc_fft_data_in_11_), 
	.A(FE_OFN1560_acc_fft_data_in_11_));
   CLKBUFX2TS FE_OFC1561_acc_fft_data_in_11_ (.Y(FE_OFN1561_acc_fft_data_in_11_), 
	.A(FE_OFN1560_acc_fft_data_in_11_));
   CLKBUFX2TS FE_OFC1560_acc_fft_data_in_11_ (.Y(FE_OFN1560_acc_fft_data_in_11_), 
	.A(FE_OFN1559_acc_fft_data_in_11_));
   CLKBUFX2TS FE_OFC1559_acc_fft_data_in_11_ (.Y(FE_OFN1559_acc_fft_data_in_11_), 
	.A(acc_fft_data_in[11]));
   CLKBUFX2TS FE_OFC1558_acc_fft_data_in_12_ (.Y(FE_OFN1558_acc_fft_data_in_12_), 
	.A(FE_OFN1557_acc_fft_data_in_12_));
   CLKBUFX2TS FE_OFC1557_acc_fft_data_in_12_ (.Y(FE_OFN1557_acc_fft_data_in_12_), 
	.A(FE_OFN1556_acc_fft_data_in_12_));
   CLKBUFX2TS FE_OFC1556_acc_fft_data_in_12_ (.Y(FE_OFN1556_acc_fft_data_in_12_), 
	.A(FE_OFN1554_acc_fft_data_in_12_));
   CLKBUFX2TS FE_OFC1555_acc_fft_data_in_12_ (.Y(FE_OFN1555_acc_fft_data_in_12_), 
	.A(FE_OFN1554_acc_fft_data_in_12_));
   CLKBUFX2TS FE_OFC1554_acc_fft_data_in_12_ (.Y(FE_OFN1554_acc_fft_data_in_12_), 
	.A(FE_OFN1553_acc_fft_data_in_12_));
   CLKBUFX2TS FE_OFC1553_acc_fft_data_in_12_ (.Y(FE_OFN1553_acc_fft_data_in_12_), 
	.A(acc_fft_data_in[12]));
   CLKBUFX2TS FE_OFC1552_acc_fft_data_in_13_ (.Y(FE_OFN1552_acc_fft_data_in_13_), 
	.A(FE_OFN1551_acc_fft_data_in_13_));
   CLKBUFX2TS FE_OFC1551_acc_fft_data_in_13_ (.Y(FE_OFN1551_acc_fft_data_in_13_), 
	.A(FE_OFN1550_acc_fft_data_in_13_));
   CLKBUFX2TS FE_OFC1550_acc_fft_data_in_13_ (.Y(FE_OFN1550_acc_fft_data_in_13_), 
	.A(FE_OFN1549_acc_fft_data_in_13_));
   CLKBUFX2TS FE_OFC1549_acc_fft_data_in_13_ (.Y(FE_OFN1549_acc_fft_data_in_13_), 
	.A(FE_OFN1548_acc_fft_data_in_13_));
   CLKBUFX2TS FE_OFC1548_acc_fft_data_in_13_ (.Y(FE_OFN1548_acc_fft_data_in_13_), 
	.A(acc_fft_data_in[13]));
   CLKBUFX2TS FE_OFC1547_acc_fft_data_in_14_ (.Y(FE_OFN1547_acc_fft_data_in_14_), 
	.A(FE_OFN1545_acc_fft_data_in_14_));
   CLKBUFX2TS FE_OFC1546_acc_fft_data_in_14_ (.Y(FE_OFN1546_acc_fft_data_in_14_), 
	.A(FE_OFN1545_acc_fft_data_in_14_));
   CLKBUFX2TS FE_OFC1545_acc_fft_data_in_14_ (.Y(FE_OFN1545_acc_fft_data_in_14_), 
	.A(FE_OFN1544_acc_fft_data_in_14_));
   CLKBUFX2TS FE_OFC1544_acc_fft_data_in_14_ (.Y(FE_OFN1544_acc_fft_data_in_14_), 
	.A(FE_OFN1543_acc_fft_data_in_14_));
   CLKBUFX2TS FE_OFC1543_acc_fft_data_in_14_ (.Y(FE_OFN1543_acc_fft_data_in_14_), 
	.A(acc_fft_data_in[14]));
   CLKBUFX2TS FE_OFC1542_acc_fft_data_in_15_ (.Y(FE_OFN1542_acc_fft_data_in_15_), 
	.A(FE_OFN1541_acc_fft_data_in_15_));
   CLKBUFX2TS FE_OFC1541_acc_fft_data_in_15_ (.Y(FE_OFN1541_acc_fft_data_in_15_), 
	.A(FE_OFN1540_acc_fft_data_in_15_));
   CLKBUFX2TS FE_OFC1540_acc_fft_data_in_15_ (.Y(FE_OFN1540_acc_fft_data_in_15_), 
	.A(FE_OFN1539_acc_fft_data_in_15_));
   CLKBUFX2TS FE_OFC1539_acc_fft_data_in_15_ (.Y(FE_OFN1539_acc_fft_data_in_15_), 
	.A(FE_OFN1538_acc_fft_data_in_15_));
   CLKBUFX2TS FE_OFC1538_acc_fft_data_in_15_ (.Y(FE_OFN1538_acc_fft_data_in_15_), 
	.A(acc_fft_data_in[15]));
   CLKBUFX2TS FE_OFC1537_acc_fft_data_in_16_ (.Y(FE_OFN1537_acc_fft_data_in_16_), 
	.A(FE_OFN1536_acc_fft_data_in_16_));
   CLKBUFX2TS FE_OFC1536_acc_fft_data_in_16_ (.Y(FE_OFN1536_acc_fft_data_in_16_), 
	.A(FE_OFN1535_acc_fft_data_in_16_));
   CLKBUFX2TS FE_OFC1535_acc_fft_data_in_16_ (.Y(FE_OFN1535_acc_fft_data_in_16_), 
	.A(FE_OFN1534_acc_fft_data_in_16_));
   CLKBUFX2TS FE_OFC1534_acc_fft_data_in_16_ (.Y(FE_OFN1534_acc_fft_data_in_16_), 
	.A(FE_OFN1533_acc_fft_data_in_16_));
   CLKBUFX2TS FE_OFC1533_acc_fft_data_in_16_ (.Y(FE_OFN1533_acc_fft_data_in_16_), 
	.A(acc_fft_data_in[16]));
   CLKBUFX2TS FE_OFC1532_acc_fft_data_in_17_ (.Y(FE_OFN1532_acc_fft_data_in_17_), 
	.A(FE_OFN1531_acc_fft_data_in_17_));
   CLKBUFX2TS FE_OFC1531_acc_fft_data_in_17_ (.Y(FE_OFN1531_acc_fft_data_in_17_), 
	.A(FE_OFN1530_acc_fft_data_in_17_));
   CLKBUFX2TS FE_OFC1530_acc_fft_data_in_17_ (.Y(FE_OFN1530_acc_fft_data_in_17_), 
	.A(FE_OFN1529_acc_fft_data_in_17_));
   CLKBUFX2TS FE_OFC1529_acc_fft_data_in_17_ (.Y(FE_OFN1529_acc_fft_data_in_17_), 
	.A(FE_OFN1528_acc_fft_data_in_17_));
   CLKBUFX2TS FE_OFC1528_acc_fft_data_in_17_ (.Y(FE_OFN1528_acc_fft_data_in_17_), 
	.A(FE_OFN1527_acc_fft_data_in_17_));
   CLKBUFX2TS FE_OFC1527_acc_fft_data_in_17_ (.Y(FE_OFN1527_acc_fft_data_in_17_), 
	.A(acc_fft_data_in[17]));
   CLKBUFX2TS FE_OFC1526_acc_fft_data_in_18_ (.Y(FE_OFN1526_acc_fft_data_in_18_), 
	.A(FE_OFN1522_acc_fft_data_in_18_));
   CLKBUFX2TS FE_OFC1525_acc_fft_data_in_18_ (.Y(FE_OFN1525_acc_fft_data_in_18_), 
	.A(FE_OFN1524_acc_fft_data_in_18_));
   CLKINVX1TS FE_OFC1524_acc_fft_data_in_18_ (.Y(FE_OFN1524_acc_fft_data_in_18_), 
	.A(FE_OFN1521_acc_fft_data_in_18_));
   CLKINVX1TS FE_OFC1523_acc_fft_data_in_18_ (.Y(FE_OFN1523_acc_fft_data_in_18_), 
	.A(FE_OFN1521_acc_fft_data_in_18_));
   CLKBUFX2TS FE_OFC1522_acc_fft_data_in_18_ (.Y(FE_OFN1522_acc_fft_data_in_18_), 
	.A(FE_OFN1520_acc_fft_data_in_18_));
   CLKINVX1TS FE_OFC1521_acc_fft_data_in_18_ (.Y(FE_OFN1521_acc_fft_data_in_18_), 
	.A(FE_OFN1520_acc_fft_data_in_18_));
   CLKBUFX2TS FE_OFC1520_acc_fft_data_in_18_ (.Y(FE_OFN1520_acc_fft_data_in_18_), 
	.A(acc_fft_data_in[18]));
   CLKBUFX2TS FE_OFC1519_acc_fft_data_in_19_ (.Y(FE_OFN1519_acc_fft_data_in_19_), 
	.A(FE_OFN1518_acc_fft_data_in_19_));
   CLKBUFX2TS FE_OFC1518_acc_fft_data_in_19_ (.Y(FE_OFN1518_acc_fft_data_in_19_), 
	.A(FE_OFN1517_acc_fft_data_in_19_));
   CLKBUFX2TS FE_OFC1517_acc_fft_data_in_19_ (.Y(FE_OFN1517_acc_fft_data_in_19_), 
	.A(FE_OFN1516_acc_fft_data_in_19_));
   CLKBUFX2TS FE_OFC1516_acc_fft_data_in_19_ (.Y(FE_OFN1516_acc_fft_data_in_19_), 
	.A(FE_OFN1515_acc_fft_data_in_19_));
   CLKBUFX2TS FE_OFC1515_acc_fft_data_in_19_ (.Y(FE_OFN1515_acc_fft_data_in_19_), 
	.A(acc_fft_data_in[19]));
   CLKBUFX2TS FE_OFC1514_acc_fft_data_in_20_ (.Y(FE_OFN1514_acc_fft_data_in_20_), 
	.A(FE_OFN1513_acc_fft_data_in_20_));
   CLKBUFX2TS FE_OFC1513_acc_fft_data_in_20_ (.Y(FE_OFN1513_acc_fft_data_in_20_), 
	.A(FE_OFN1512_acc_fft_data_in_20_));
   CLKBUFX2TS FE_OFC1512_acc_fft_data_in_20_ (.Y(FE_OFN1512_acc_fft_data_in_20_), 
	.A(FE_OFN1511_acc_fft_data_in_20_));
   CLKBUFX2TS FE_OFC1511_acc_fft_data_in_20_ (.Y(FE_OFN1511_acc_fft_data_in_20_), 
	.A(FE_OFN1510_acc_fft_data_in_20_));
   CLKBUFX2TS FE_OFC1510_acc_fft_data_in_20_ (.Y(FE_OFN1510_acc_fft_data_in_20_), 
	.A(acc_fft_data_in[20]));
   CLKBUFX2TS FE_OFC1509_acc_fft_data_in_21_ (.Y(FE_OFN1509_acc_fft_data_in_21_), 
	.A(FE_OFN1507_acc_fft_data_in_21_));
   CLKBUFX2TS FE_OFC1508_acc_fft_data_in_21_ (.Y(FE_OFN1508_acc_fft_data_in_21_), 
	.A(FE_OFN1506_acc_fft_data_in_21_));
   CLKBUFX2TS FE_OFC1507_acc_fft_data_in_21_ (.Y(FE_OFN1507_acc_fft_data_in_21_), 
	.A(FE_OFN1505_acc_fft_data_in_21_));
   CLKBUFX2TS FE_OFC1506_acc_fft_data_in_21_ (.Y(FE_OFN1506_acc_fft_data_in_21_), 
	.A(FE_OFN1505_acc_fft_data_in_21_));
   CLKBUFX2TS FE_OFC1505_acc_fft_data_in_21_ (.Y(FE_OFN1505_acc_fft_data_in_21_), 
	.A(acc_fft_data_in[21]));
   CLKINVX1TS FE_OFC1504_acc_fft_data_in_22_ (.Y(FE_OFN1504_acc_fft_data_in_22_), 
	.A(FE_OFN1502_acc_fft_data_in_22_));
   CLKINVX1TS FE_OFC1503_acc_fft_data_in_22_ (.Y(FE_OFN1503_acc_fft_data_in_22_), 
	.A(FE_OFN1502_acc_fft_data_in_22_));
   CLKINVX1TS FE_OFC1502_acc_fft_data_in_22_ (.Y(FE_OFN1502_acc_fft_data_in_22_), 
	.A(FE_OFN1499_acc_fft_data_in_22_));
   CLKBUFX2TS FE_OFC1501_acc_fft_data_in_22_ (.Y(FE_OFN1501_acc_fft_data_in_22_), 
	.A(FE_OFN1500_acc_fft_data_in_22_));
   CLKBUFX2TS FE_OFC1500_acc_fft_data_in_22_ (.Y(FE_OFN1500_acc_fft_data_in_22_), 
	.A(FE_OFN1499_acc_fft_data_in_22_));
   CLKBUFX2TS FE_OFC1499_acc_fft_data_in_22_ (.Y(FE_OFN1499_acc_fft_data_in_22_), 
	.A(FE_OFN1498_acc_fft_data_in_22_));
   CLKBUFX2TS FE_OFC1498_acc_fft_data_in_22_ (.Y(FE_OFN1498_acc_fft_data_in_22_), 
	.A(acc_fft_data_in[22]));
   CLKBUFX2TS FE_OFC1497_acc_fft_data_in_23_ (.Y(FE_OFN1497_acc_fft_data_in_23_), 
	.A(FE_OFN1496_acc_fft_data_in_23_));
   CLKBUFX2TS FE_OFC1496_acc_fft_data_in_23_ (.Y(FE_OFN1496_acc_fft_data_in_23_), 
	.A(FE_OFN1493_acc_fft_data_in_23_));
   CLKBUFX2TS FE_OFC1495_acc_fft_data_in_23_ (.Y(FE_OFN1495_acc_fft_data_in_23_), 
	.A(FE_OFN1493_acc_fft_data_in_23_));
   CLKBUFX2TS FE_OFC1494_acc_fft_data_in_23_ (.Y(FE_OFN1494_acc_fft_data_in_23_), 
	.A(FE_OFN1493_acc_fft_data_in_23_));
   CLKBUFX2TS FE_OFC1493_acc_fft_data_in_23_ (.Y(FE_OFN1493_acc_fft_data_in_23_), 
	.A(acc_fft_data_in[23]));
   CLKBUFX2TS FE_OFC1492_acc_fft_data_in_24_ (.Y(FE_OFN1492_acc_fft_data_in_24_), 
	.A(FE_OFN1489_acc_fft_data_in_24_));
   CLKBUFX2TS FE_OFC1491_acc_fft_data_in_24_ (.Y(FE_OFN1491_acc_fft_data_in_24_), 
	.A(FE_OFN1490_acc_fft_data_in_24_));
   CLKBUFX2TS FE_OFC1490_acc_fft_data_in_24_ (.Y(FE_OFN1490_acc_fft_data_in_24_), 
	.A(FE_OFN1488_acc_fft_data_in_24_));
   CLKBUFX2TS FE_OFC1489_acc_fft_data_in_24_ (.Y(FE_OFN1489_acc_fft_data_in_24_), 
	.A(FE_OFN1488_acc_fft_data_in_24_));
   CLKBUFX2TS FE_OFC1488_acc_fft_data_in_24_ (.Y(FE_OFN1488_acc_fft_data_in_24_), 
	.A(acc_fft_data_in[24]));
   CLKBUFX2TS FE_OFC1487_acc_fft_data_in_25_ (.Y(FE_OFN1487_acc_fft_data_in_25_), 
	.A(FE_OFN1485_acc_fft_data_in_25_));
   CLKBUFX2TS FE_OFC1486_acc_fft_data_in_25_ (.Y(FE_OFN1486_acc_fft_data_in_25_), 
	.A(FE_OFN1484_acc_fft_data_in_25_));
   CLKBUFX2TS FE_OFC1485_acc_fft_data_in_25_ (.Y(FE_OFN1485_acc_fft_data_in_25_), 
	.A(FE_OFN1484_acc_fft_data_in_25_));
   CLKBUFX2TS FE_OFC1484_acc_fft_data_in_25_ (.Y(FE_OFN1484_acc_fft_data_in_25_), 
	.A(FE_OFN1483_acc_fft_data_in_25_));
   CLKBUFX2TS FE_OFC1483_acc_fft_data_in_25_ (.Y(FE_OFN1483_acc_fft_data_in_25_), 
	.A(acc_fft_data_in[25]));
   CLKBUFX2TS FE_OFC1482_acc_fft_data_in_26_ (.Y(FE_OFN1482_acc_fft_data_in_26_), 
	.A(FE_OFN1481_acc_fft_data_in_26_));
   CLKBUFX2TS FE_OFC1481_acc_fft_data_in_26_ (.Y(FE_OFN1481_acc_fft_data_in_26_), 
	.A(FE_OFN1480_acc_fft_data_in_26_));
   CLKBUFX2TS FE_OFC1480_acc_fft_data_in_26_ (.Y(FE_OFN1480_acc_fft_data_in_26_), 
	.A(FE_OFN1479_acc_fft_data_in_26_));
   CLKBUFX2TS FE_OFC1479_acc_fft_data_in_26_ (.Y(FE_OFN1479_acc_fft_data_in_26_), 
	.A(FE_OFN1478_acc_fft_data_in_26_));
   CLKBUFX2TS FE_OFC1478_acc_fft_data_in_26_ (.Y(FE_OFN1478_acc_fft_data_in_26_), 
	.A(acc_fft_data_in[26]));
   CLKBUFX2TS FE_OFC1477_acc_fft_data_in_27_ (.Y(FE_OFN1477_acc_fft_data_in_27_), 
	.A(FE_OFN1476_acc_fft_data_in_27_));
   CLKBUFX2TS FE_OFC1476_acc_fft_data_in_27_ (.Y(FE_OFN1476_acc_fft_data_in_27_), 
	.A(FE_OFN1475_acc_fft_data_in_27_));
   CLKBUFX2TS FE_OFC1475_acc_fft_data_in_27_ (.Y(FE_OFN1475_acc_fft_data_in_27_), 
	.A(FE_OFN1474_acc_fft_data_in_27_));
   CLKBUFX2TS FE_OFC1474_acc_fft_data_in_27_ (.Y(FE_OFN1474_acc_fft_data_in_27_), 
	.A(FE_OFN1473_acc_fft_data_in_27_));
   CLKBUFX2TS FE_OFC1473_acc_fft_data_in_27_ (.Y(FE_OFN1473_acc_fft_data_in_27_), 
	.A(acc_fft_data_in[27]));
   CLKBUFX2TS FE_OFC1472_acc_fft_data_in_28_ (.Y(FE_OFN1472_acc_fft_data_in_28_), 
	.A(FE_OFN1470_acc_fft_data_in_28_));
   CLKBUFX2TS FE_OFC1471_acc_fft_data_in_28_ (.Y(FE_OFN1471_acc_fft_data_in_28_), 
	.A(FE_OFN1820_acc_fft_data_in_28_));
   CLKBUFX2TS FE_OFC1470_acc_fft_data_in_28_ (.Y(FE_OFN1470_acc_fft_data_in_28_), 
	.A(FE_OFN1821_acc_fft_data_in_28_));
   CLKBUFX2TS FE_OFC1469_acc_fft_data_in_28_ (.Y(FE_OFN1469_acc_fft_data_in_28_), 
	.A(FE_OFN1468_acc_fft_data_in_28_));
   CLKBUFX2TS FE_OFC1468_acc_fft_data_in_28_ (.Y(FE_OFN1468_acc_fft_data_in_28_), 
	.A(acc_fft_data_in[28]));
   CLKBUFX2TS FE_OFC1467_acc_fft_data_in_29_ (.Y(FE_OFN1467_acc_fft_data_in_29_), 
	.A(FE_OFN1465_acc_fft_data_in_29_));
   CLKBUFX2TS FE_OFC1466_acc_fft_data_in_29_ (.Y(FE_OFN1466_acc_fft_data_in_29_), 
	.A(FE_OFN1464_acc_fft_data_in_29_));
   CLKBUFX2TS FE_OFC1465_acc_fft_data_in_29_ (.Y(FE_OFN1465_acc_fft_data_in_29_), 
	.A(FE_OFN1463_acc_fft_data_in_29_));
   CLKBUFX2TS FE_OFC1464_acc_fft_data_in_29_ (.Y(FE_OFN1464_acc_fft_data_in_29_), 
	.A(FE_OFN1463_acc_fft_data_in_29_));
   CLKBUFX2TS FE_OFC1463_acc_fft_data_in_29_ (.Y(FE_OFN1463_acc_fft_data_in_29_), 
	.A(acc_fft_data_in[29]));
   CLKBUFX2TS FE_OFC1462_acc_fft_data_in_30_ (.Y(FE_OFN1462_acc_fft_data_in_30_), 
	.A(FE_OFN1459_acc_fft_data_in_30_));
   CLKBUFX2TS FE_OFC1461_acc_fft_data_in_30_ (.Y(FE_OFN1461_acc_fft_data_in_30_), 
	.A(FE_OFN1460_acc_fft_data_in_30_));
   CLKBUFX2TS FE_OFC1460_acc_fft_data_in_30_ (.Y(FE_OFN1460_acc_fft_data_in_30_), 
	.A(FE_OFN1458_acc_fft_data_in_30_));
   CLKBUFX2TS FE_OFC1459_acc_fft_data_in_30_ (.Y(FE_OFN1459_acc_fft_data_in_30_), 
	.A(FE_OFN1458_acc_fft_data_in_30_));
   CLKBUFX2TS FE_OFC1458_acc_fft_data_in_30_ (.Y(FE_OFN1458_acc_fft_data_in_30_), 
	.A(acc_fft_data_in[30]));
   CLKBUFX2TS FE_OFC1457_acc_fft_data_in_31_ (.Y(FE_OFN1457_acc_fft_data_in_31_), 
	.A(FE_OFN1455_acc_fft_data_in_31_));
   CLKBUFX2TS FE_OFC1456_acc_fft_data_in_31_ (.Y(FE_OFN1456_acc_fft_data_in_31_), 
	.A(FE_OFN1454_acc_fft_data_in_31_));
   CLKBUFX2TS FE_OFC1455_acc_fft_data_in_31_ (.Y(FE_OFN1455_acc_fft_data_in_31_), 
	.A(FE_OFN1452_acc_fft_data_in_31_));
   CLKBUFX2TS FE_OFC1454_acc_fft_data_in_31_ (.Y(FE_OFN1454_acc_fft_data_in_31_), 
	.A(FE_OFN1452_acc_fft_data_in_31_));
   CLKBUFX2TS FE_OFC1453_acc_fft_data_in_31_ (.Y(FE_OFN1453_acc_fft_data_in_31_), 
	.A(FE_OFN1452_acc_fft_data_in_31_));
   CLKBUFX2TS FE_OFC1452_acc_fft_data_in_31_ (.Y(FE_OFN1452_acc_fft_data_in_31_), 
	.A(acc_fft_data_in[31]));
   CLKBUFX2TS FE_OFC1451_acc_fir_put (.Y(FE_OFN1451_acc_fir_put), 
	.A(acc_fir_put));
   CLKBUFX2TS FE_OFC1450_acc_fir_get (.Y(FE_OFN1450_acc_fir_get), 
	.A(acc_fir_get));
   CLKBUFX2TS FE_OFC1449_acc_fft_put (.Y(FE_OFN1449_acc_fft_put), 
	.A(acc_fft_put));
   CLKBUFX2TS FE_OFC1448_acc_fft_get (.Y(FE_OFN1448_acc_fft_get), 
	.A(acc_fft_get));
   CLKBUFX2TS FE_OFC1447_reset (.Y(FE_OFN1447_reset), 
	.A(reset));
   CLKBUFX2TS FE_OFC1446_router_addr_calc_fir_read_calc_count_0_ (.Y(FE_OFN1446_router_addr_calc_fir_read_calc_count_0_), 
	.A(\router/addr_calc/fir_read_calc/count[0] ));
   CLKBUFX2TS FE_OFC1445_router_addr_calc_fir_write_calc_count_0_ (.Y(FE_OFN1445_router_addr_calc_fir_write_calc_count_0_), 
	.A(\router/addr_calc/fir_write_calc/count[0] ));
   CLKBUFX2TS FE_OFC1444_router_addr_calc_fft_read_calc_count_0_ (.Y(FE_OFN1444_router_addr_calc_fft_read_calc_count_0_), 
	.A(\router/addr_calc/fft_read_calc/count[0] ));
   CLKBUFX2TS FE_OFC1443_router_addr_calc_fft_write_calc_count_0_ (.Y(FE_OFN1443_router_addr_calc_fft_write_calc_count_0_), 
	.A(\router/addr_calc/fft_write_calc/count[0] ));
   CLKBUFX2TS FE_OFC1442_router_addr_calc_iir_write_calc_count_0_ (.Y(FE_OFN1442_router_addr_calc_iir_write_calc_count_0_), 
	.A(\router/addr_calc/iir_write_calc/count[0] ));
   CLKBUFX2TS FE_OFC1441_router_addr_calc_iir_write_calc_count_16_ (.Y(FE_OFN1441_router_addr_calc_iir_write_calc_count_16_), 
	.A(\router/addr_calc/iir_write_calc/count[16] ));
   CLKBUFX2TS FE_OFC1440_router_addr_calc_iir_write_calc_count_19_ (.Y(FE_OFN1440_router_addr_calc_iir_write_calc_count_19_), 
	.A(\router/addr_calc/iir_write_calc/count[19] ));
   CLKBUFX2TS FE_OFC1439_router_addr_calc_iir_write_calc_count_27_ (.Y(FE_OFN1439_router_addr_calc_iir_write_calc_count_27_), 
	.A(\router/addr_calc/iir_write_calc/count[27] ));
   CLKBUFX2TS FE_OFC1438_router_data_from_fft (.Y(FE_OFN1438_router_data_from_fft), 
	.A(\router/data_from_fft ));
   CLKBUFX2TS FE_OFC1437_n8093 (.Y(FE_OFN1437_n8093), 
	.A(FE_OFN1436_n8093));
   CLKBUFX2TS FE_OFC1436_n8093 (.Y(FE_OFN1436_n8093), 
	.A(FE_OFN1434_n8093));
   CLKBUFX2TS FE_OFC1435_n8093 (.Y(FE_OFN1435_n8093), 
	.A(FE_OFN1434_n8093));
   CLKBUFX2TS FE_OFC1434_n8093 (.Y(FE_OFN1434_n8093), 
	.A(FE_OFN1433_n8093));
   CLKBUFX2TS FE_OFC1433_n8093 (.Y(FE_OFN1433_n8093), 
	.A(n8093));
   CLKBUFX2TS FE_OFC1432_n8092 (.Y(FE_OFN1432_n8092), 
	.A(FE_OFN1430_n8092));
   CLKBUFX2TS FE_OFC1431_n8092 (.Y(FE_OFN1431_n8092), 
	.A(n8092));
   CLKBUFX2TS FE_OFC1430_n8092 (.Y(FE_OFN1430_n8092), 
	.A(FE_OFN1429_n8092));
   CLKBUFX2TS FE_OFC1429_n8092 (.Y(FE_OFN1429_n8092), 
	.A(n8092));
   CLKBUFX2TS FE_OFC1428_n8091 (.Y(FE_OFN1428_n8091), 
	.A(FE_OFN1425_n8091));
   CLKBUFX2TS FE_OFC1427_n8091 (.Y(FE_OFN1427_n8091), 
	.A(FE_OFN1425_n8091));
   CLKBUFX2TS FE_OFC1426_n8091 (.Y(FE_OFN1426_n8091), 
	.A(n8091));
   CLKBUFX2TS FE_OFC1425_n8091 (.Y(FE_OFN1425_n8091), 
	.A(n8091));
   CLKBUFX2TS FE_OFC1424_n8090 (.Y(FE_OFN1424_n8090), 
	.A(FE_OFN1422_n8090));
   CLKBUFX2TS FE_OFC1423_n8090 (.Y(FE_OFN1423_n8090), 
	.A(FE_OFN1422_n8090));
   CLKBUFX2TS FE_OFC1422_n8090 (.Y(FE_OFN1422_n8090), 
	.A(FE_OFN1420_n8090));
   CLKBUFX2TS FE_OFC1421_n8090 (.Y(FE_OFN1421_n8090), 
	.A(FE_OFN1420_n8090));
   CLKBUFX2TS FE_OFC1420_n8090 (.Y(FE_OFN1420_n8090), 
	.A(n8090));
   CLKBUFX2TS FE_OFC1419_n8089 (.Y(FE_OFN1419_n8089), 
	.A(FE_OFN1417_n8089));
   CLKBUFX2TS FE_OFC1418_n8089 (.Y(FE_OFN1418_n8089), 
	.A(FE_OFN1417_n8089));
   CLKBUFX2TS FE_OFC1417_n8089 (.Y(FE_OFN1417_n8089), 
	.A(FE_OFN1416_n8089));
   CLKBUFX2TS FE_OFC1416_n8089 (.Y(FE_OFN1416_n8089), 
	.A(n8089));
   CLKBUFX2TS FE_OFC1415_n8088 (.Y(FE_OFN1415_n8088), 
	.A(FE_OFN1414_n8088));
   CLKBUFX2TS FE_OFC1414_n8088 (.Y(FE_OFN1414_n8088), 
	.A(FE_OFN1413_n8088));
   CLKBUFX2TS FE_OFC1413_n8088 (.Y(FE_OFN1413_n8088), 
	.A(FE_OFN1412_n8088));
   CLKBUFX2TS FE_OFC1412_n8088 (.Y(FE_OFN1412_n8088), 
	.A(n8088));
   CLKBUFX2TS FE_OFC1411_n8087 (.Y(FE_OFN1411_n8087), 
	.A(FE_OFN1409_n8087));
   CLKBUFX2TS FE_OFC1410_n8087 (.Y(FE_OFN1410_n8087), 
	.A(FE_OFN1409_n8087));
   CLKBUFX2TS FE_OFC1409_n8087 (.Y(FE_OFN1409_n8087), 
	.A(FE_OFN1408_n8087));
   CLKBUFX2TS FE_OFC1408_n8087 (.Y(FE_OFN1408_n8087), 
	.A(FE_OFN1407_n8087));
   CLKBUFX2TS FE_OFC1407_n8087 (.Y(FE_OFN1407_n8087), 
	.A(n8087));
   CLKBUFX2TS FE_OFC1406_n8086 (.Y(FE_OFN1406_n8086), 
	.A(FE_OFN1404_n8086));
   CLKBUFX2TS FE_OFC1405_n8086 (.Y(FE_OFN1405_n8086), 
	.A(FE_OFN1404_n8086));
   CLKBUFX2TS FE_OFC1404_n8086 (.Y(FE_OFN1404_n8086), 
	.A(FE_OFN1403_n8086));
   CLKBUFX2TS FE_OFC1403_n8086 (.Y(FE_OFN1403_n8086), 
	.A(n8086));
   CLKBUFX2TS FE_OFC1402_n8085 (.Y(FE_OFN1402_n8085), 
	.A(FE_OFN1401_n8085));
   CLKBUFX2TS FE_OFC1401_n8085 (.Y(FE_OFN1401_n8085), 
	.A(FE_OFN1400_n8085));
   CLKBUFX2TS FE_OFC1400_n8085 (.Y(FE_OFN1400_n8085), 
	.A(FE_OFN1399_n8085));
   CLKBUFX2TS FE_OFC1399_n8085 (.Y(FE_OFN1399_n8085), 
	.A(n8085));
   CLKBUFX2TS FE_OFC1398_n8084 (.Y(FE_OFN1398_n8084), 
	.A(FE_OFN1397_n8084));
   CLKBUFX2TS FE_OFC1397_n8084 (.Y(FE_OFN1397_n8084), 
	.A(FE_OFN1396_n8084));
   CLKBUFX2TS FE_OFC1396_n8084 (.Y(FE_OFN1396_n8084), 
	.A(FE_OFN1395_n8084));
   CLKBUFX2TS FE_OFC1395_n8084 (.Y(FE_OFN1395_n8084), 
	.A(FE_OFN1394_n8084));
   CLKBUFX2TS FE_OFC1394_n8084 (.Y(FE_OFN1394_n8084), 
	.A(n8084));
   CLKBUFX2TS FE_OFC1393_n8083 (.Y(FE_OFN1393_n8083), 
	.A(FE_OFN1391_n8083));
   CLKBUFX2TS FE_OFC1392_n8083 (.Y(FE_OFN1392_n8083), 
	.A(FE_OFN1391_n8083));
   CLKBUFX2TS FE_OFC1391_n8083 (.Y(FE_OFN1391_n8083), 
	.A(FE_OFN1390_n8083));
   CLKBUFX2TS FE_OFC1390_n8083 (.Y(FE_OFN1390_n8083), 
	.A(n8083));
   CLKBUFX2TS FE_OFC1389_n8083 (.Y(FE_OFN1389_n8083), 
	.A(n8083));
   CLKBUFX2TS FE_OFC1388_n8082 (.Y(FE_OFN1388_n8082), 
	.A(FE_OFN1387_n8082));
   CLKBUFX2TS FE_OFC1387_n8082 (.Y(FE_OFN1387_n8082), 
	.A(FE_OFN1385_n8082));
   CLKBUFX2TS FE_OFC1386_n8082 (.Y(FE_OFN1386_n8082), 
	.A(FE_OFN1384_n8082));
   CLKBUFX2TS FE_OFC1385_n8082 (.Y(FE_OFN1385_n8082), 
	.A(n8082));
   CLKBUFX2TS FE_OFC1384_n8082 (.Y(FE_OFN1384_n8082), 
	.A(n8082));
   CLKBUFX2TS FE_OFC1383_n8081 (.Y(FE_OFN1383_n8081), 
	.A(FE_OFN1381_n8081));
   CLKBUFX2TS FE_OFC1382_n8081 (.Y(FE_OFN1382_n8081), 
	.A(FE_OFN1380_n8081));
   CLKBUFX2TS FE_OFC1381_n8081 (.Y(FE_OFN1381_n8081), 
	.A(n8081));
   CLKBUFX2TS FE_OFC1380_n8081 (.Y(FE_OFN1380_n8081), 
	.A(n8081));
   CLKBUFX2TS FE_OFC1379_n8080 (.Y(FE_OFN1379_n8080), 
	.A(FE_OFN1378_n8080));
   CLKBUFX2TS FE_OFC1378_n8080 (.Y(FE_OFN1378_n8080), 
	.A(FE_OFN1376_n8080));
   CLKBUFX2TS FE_OFC1377_n8080 (.Y(FE_OFN1377_n8080), 
	.A(n8080));
   CLKBUFX2TS FE_OFC1376_n8080 (.Y(FE_OFN1376_n8080), 
	.A(n8080));
   CLKBUFX2TS FE_OFC1375_n8078 (.Y(FE_OFN1375_n8078), 
	.A(FE_OFN1374_n8078));
   CLKBUFX2TS FE_OFC1374_n8078 (.Y(FE_OFN1374_n8078), 
	.A(FE_OFN1373_n8078));
   CLKBUFX2TS FE_OFC1373_n8078 (.Y(FE_OFN1373_n8078), 
	.A(FE_OFN1372_n8078));
   CLKBUFX2TS FE_OFC1372_n8078 (.Y(FE_OFN1372_n8078), 
	.A(FE_OFN1371_n8078));
   CLKBUFX2TS FE_OFC1371_n8078 (.Y(FE_OFN1371_n8078), 
	.A(n8078));
   CLKBUFX2TS FE_OFC1370_n8077 (.Y(FE_OFN1370_n8077), 
	.A(FE_OFN1369_n8077));
   CLKBUFX2TS FE_OFC1369_n8077 (.Y(FE_OFN1369_n8077), 
	.A(FE_OFN1367_n8077));
   CLKBUFX2TS FE_OFC1368_n8077 (.Y(FE_OFN1368_n8077), 
	.A(FE_OFN1367_n8077));
   CLKBUFX2TS FE_OFC1367_n8077 (.Y(FE_OFN1367_n8077), 
	.A(FE_OFN1366_n8077));
   CLKBUFX2TS FE_OFC1366_n8077 (.Y(FE_OFN1366_n8077), 
	.A(n8077));
   CLKBUFX2TS FE_OFC1365_n8076 (.Y(FE_OFN1365_n8076), 
	.A(FE_OFN1364_n8076));
   CLKBUFX2TS FE_OFC1364_n8076 (.Y(FE_OFN1364_n8076), 
	.A(FE_OFN1363_n8076));
   CLKBUFX2TS FE_OFC1363_n8076 (.Y(FE_OFN1363_n8076), 
	.A(FE_OFN1362_n8076));
   CLKBUFX2TS FE_OFC1362_n8076 (.Y(FE_OFN1362_n8076), 
	.A(n8076));
   CLKBUFX2TS FE_OFC1361_n8075 (.Y(FE_OFN1361_n8075), 
	.A(FE_OFN1360_n8075));
   CLKBUFX2TS FE_OFC1360_n8075 (.Y(FE_OFN1360_n8075), 
	.A(FE_OFN1358_n8075));
   CLKBUFX2TS FE_OFC1359_n8075 (.Y(FE_OFN1359_n8075), 
	.A(FE_OFN1358_n8075));
   CLKBUFX2TS FE_OFC1358_n8075 (.Y(FE_OFN1358_n8075), 
	.A(FE_OFN1357_n8075));
   CLKBUFX2TS FE_OFC1357_n8075 (.Y(FE_OFN1357_n8075), 
	.A(n8075));
   CLKBUFX2TS FE_OFC1356_n8074 (.Y(FE_OFN1356_n8074), 
	.A(FE_OFN1355_n8074));
   CLKBUFX2TS FE_OFC1355_n8074 (.Y(FE_OFN1355_n8074), 
	.A(FE_OFN1354_n8074));
   CLKBUFX2TS FE_OFC1354_n8074 (.Y(FE_OFN1354_n8074), 
	.A(FE_OFN1353_n8074));
   CLKBUFX2TS FE_OFC1353_n8074 (.Y(FE_OFN1353_n8074), 
	.A(n8074));
   CLKBUFX2TS FE_OFC1352_n8073 (.Y(FE_OFN1352_n8073), 
	.A(FE_OFN1351_n8073));
   CLKBUFX2TS FE_OFC1351_n8073 (.Y(FE_OFN1351_n8073), 
	.A(FE_OFN1350_n8073));
   CLKBUFX2TS FE_OFC1350_n8073 (.Y(FE_OFN1350_n8073), 
	.A(n8073));
   CLKBUFX2TS FE_OFC1349_n8073 (.Y(FE_OFN1349_n8073), 
	.A(n8073));
   CLKBUFX2TS FE_OFC1348_n8072 (.Y(FE_OFN1348_n8072), 
	.A(FE_OFN1347_n8072));
   CLKBUFX2TS FE_OFC1347_n8072 (.Y(FE_OFN1347_n8072), 
	.A(FE_OFN1345_n8072));
   CLKBUFX2TS FE_OFC1346_n8072 (.Y(FE_OFN1346_n8072), 
	.A(FE_OFN1345_n8072));
   CLKBUFX2TS FE_OFC1345_n8072 (.Y(FE_OFN1345_n8072), 
	.A(FE_OFN1344_n8072));
   CLKBUFX2TS FE_OFC1344_n8072 (.Y(FE_OFN1344_n8072), 
	.A(n8072));
   CLKBUFX2TS FE_OFC1343_n8071 (.Y(FE_OFN1343_n8071), 
	.A(FE_OFN1342_n8071));
   CLKBUFX2TS FE_OFC1342_n8071 (.Y(FE_OFN1342_n8071), 
	.A(FE_OFN1341_n8071));
   CLKBUFX2TS FE_OFC1341_n8071 (.Y(FE_OFN1341_n8071), 
	.A(FE_OFN1340_n8071));
   CLKBUFX2TS FE_OFC1340_n8071 (.Y(FE_OFN1340_n8071), 
	.A(FE_OFN1339_n8071));
   CLKBUFX2TS FE_OFC1339_n8071 (.Y(FE_OFN1339_n8071), 
	.A(n8071));
   CLKBUFX2TS FE_OFC1338_n8070 (.Y(FE_OFN1338_n8070), 
	.A(FE_OFN1337_n8070));
   CLKBUFX2TS FE_OFC1337_n8070 (.Y(FE_OFN1337_n8070), 
	.A(FE_OFN1336_n8070));
   CLKBUFX2TS FE_OFC1336_n8070 (.Y(FE_OFN1336_n8070), 
	.A(FE_OFN1335_n8070));
   CLKBUFX2TS FE_OFC1335_n8070 (.Y(FE_OFN1335_n8070), 
	.A(n8070));
   CLKBUFX2TS FE_OFC1334_n8069 (.Y(FE_OFN1334_n8069), 
	.A(FE_OFN1333_n8069));
   CLKBUFX2TS FE_OFC1333_n8069 (.Y(FE_OFN1333_n8069), 
	.A(FE_OFN1332_n8069));
   CLKBUFX2TS FE_OFC1332_n8069 (.Y(FE_OFN1332_n8069), 
	.A(FE_OFN1331_n8069));
   CLKBUFX2TS FE_OFC1331_n8069 (.Y(FE_OFN1331_n8069), 
	.A(n8069));
   CLKBUFX2TS FE_OFC1330_n8068 (.Y(FE_OFN1330_n8068), 
	.A(FE_OFN1329_n8068));
   CLKBUFX2TS FE_OFC1329_n8068 (.Y(FE_OFN1329_n8068), 
	.A(FE_OFN1328_n8068));
   CLKBUFX2TS FE_OFC1328_n8068 (.Y(FE_OFN1328_n8068), 
	.A(FE_OFN1327_n8068));
   CLKBUFX2TS FE_OFC1327_n8068 (.Y(FE_OFN1327_n8068), 
	.A(n8068));
   CLKBUFX2TS FE_OFC1326_n8067 (.Y(FE_OFN1326_n8067), 
	.A(FE_OFN1324_n8067));
   CLKBUFX2TS FE_OFC1325_n8067 (.Y(FE_OFN1325_n8067), 
	.A(FE_OFN1324_n8067));
   CLKBUFX2TS FE_OFC1324_n8067 (.Y(FE_OFN1324_n8067), 
	.A(FE_OFN1323_n8067));
   CLKBUFX2TS FE_OFC1323_n8067 (.Y(FE_OFN1323_n8067), 
	.A(n8067));
   CLKBUFX2TS FE_OFC1322_n8066 (.Y(FE_OFN1322_n8066), 
	.A(FE_OFN1321_n8066));
   CLKBUFX2TS FE_OFC1321_n8066 (.Y(FE_OFN1321_n8066), 
	.A(FE_OFN1320_n8066));
   CLKBUFX2TS FE_OFC1320_n8066 (.Y(FE_OFN1320_n8066), 
	.A(FE_OFN1319_n8066));
   CLKBUFX2TS FE_OFC1319_n8066 (.Y(FE_OFN1319_n8066), 
	.A(FE_OFN1318_n8066));
   CLKBUFX2TS FE_OFC1318_n8066 (.Y(FE_OFN1318_n8066), 
	.A(n8066));
   CLKBUFX2TS FE_OFC1317_n8065 (.Y(FE_OFN1317_n8065), 
	.A(FE_OFN1316_n8065));
   CLKBUFX2TS FE_OFC1316_n8065 (.Y(FE_OFN1316_n8065), 
	.A(FE_OFN1315_n8065));
   CLKBUFX2TS FE_OFC1315_n8065 (.Y(FE_OFN1315_n8065), 
	.A(FE_OFN1314_n8065));
   CLKBUFX2TS FE_OFC1314_n8065 (.Y(FE_OFN1314_n8065), 
	.A(n8065));
   CLKBUFX2TS FE_OFC1313_n8094 (.Y(FE_OFN1313_n8094), 
	.A(FE_OFN1310_n8094));
   CLKBUFX2TS FE_OFC1312_n8094 (.Y(FE_OFN1312_n8094), 
	.A(FE_OFN1311_n8094));
   CLKBUFX2TS FE_OFC1311_n8094 (.Y(FE_OFN1311_n8094), 
	.A(n8094));
   CLKBUFX2TS FE_OFC1310_n8094 (.Y(FE_OFN1310_n8094), 
	.A(n8094));
   CLKBUFX2TS FE_OFC1309_n8079 (.Y(FE_OFN1309_n8079), 
	.A(FE_OFN1308_n8079));
   CLKBUFX2TS FE_OFC1308_n8079 (.Y(FE_OFN1308_n8079), 
	.A(FE_OFN1307_n8079));
   CLKBUFX2TS FE_OFC1307_n8079 (.Y(FE_OFN1307_n8079), 
	.A(FE_OFN1306_n8079));
   CLKBUFX2TS FE_OFC1306_n8079 (.Y(FE_OFN1306_n8079), 
	.A(n8079));
   CLKBUFX2TS FE_OFC1305_n8060 (.Y(FE_OFN1305_n8060), 
	.A(FE_OFN1304_n8060));
   CLKBUFX2TS FE_OFC1304_n8060 (.Y(FE_OFN1304_n8060), 
	.A(FE_OFN1302_n8060));
   CLKBUFX2TS FE_OFC1303_n8060 (.Y(FE_OFN1303_n8060), 
	.A(FE_OFN1302_n8060));
   CLKBUFX2TS FE_OFC1302_n8060 (.Y(FE_OFN1302_n8060), 
	.A(FE_OFN1301_n8060));
   CLKBUFX2TS FE_OFC1301_n8060 (.Y(FE_OFN1301_n8060), 
	.A(n8060));
   CLKBUFX2TS FE_OFC1300_iir_enable (.Y(FE_OFN1300_iir_enable), 
	.A(FE_OFN1299_iir_enable));
   CLKBUFX2TS FE_OFC1299_iir_enable (.Y(FE_OFN1299_iir_enable), 
	.A(FE_OFN1298_iir_enable));
   CLKBUFX2TS FE_OFC1298_iir_enable (.Y(FE_OFN1298_iir_enable), 
	.A(FE_OFN1294_iir_enable));
   CLKBUFX2TS FE_OFC1297_iir_enable (.Y(FE_OFN1297_iir_enable), 
	.A(FE_OFN1294_iir_enable));
   CLKBUFX2TS FE_OFC1296_iir_enable (.Y(FE_OFN1296_iir_enable), 
	.A(FE_OFN1293_iir_enable));
   CLKBUFX2TS FE_OFC1295_iir_enable (.Y(FE_OFN1295_iir_enable), 
	.A(FE_OFN1293_iir_enable));
   CLKBUFX2TS FE_OFC1294_iir_enable (.Y(FE_OFN1294_iir_enable), 
	.A(FE_OFN1292_iir_enable));
   CLKBUFX2TS FE_OFC1293_iir_enable (.Y(FE_OFN1293_iir_enable), 
	.A(FE_OFN1291_iir_enable));
   CLKBUFX2TS FE_OFC1292_iir_enable (.Y(FE_OFN1292_iir_enable), 
	.A(FE_OFN1290_iir_enable));
   CLKBUFX2TS FE_OFC1291_iir_enable (.Y(FE_OFN1291_iir_enable), 
	.A(FE_OFN1290_iir_enable));
   CLKBUFX2TS FE_OFC1290_iir_enable (.Y(FE_OFN1290_iir_enable), 
	.A(FE_OFN1288_iir_enable));
   CLKBUFX2TS FE_OFC1289_iir_enable (.Y(FE_OFN1289_iir_enable), 
	.A(FE_OFN1288_iir_enable));
   CLKBUFX2TS FE_OFC1288_iir_enable (.Y(FE_OFN1288_iir_enable), 
	.A(FE_OFN1287_iir_enable));
   CLKBUFX2TS FE_OFC1287_iir_enable (.Y(FE_OFN1287_iir_enable), 
	.A(FE_OFN1286_iir_enable));
   CLKBUFX2TS FE_OFC1286_iir_enable (.Y(FE_OFN1286_iir_enable), 
	.A(iir_enable));
   CLKBUFX2TS FE_OFC1285_router_ram_read_enable_reg (.Y(FE_OFN1285_router_ram_read_enable_reg), 
	.A(FE_OFN1284_router_ram_read_enable_reg));
   CLKBUFX2TS FE_OFC1284_router_ram_read_enable_reg (.Y(FE_OFN1284_router_ram_read_enable_reg), 
	.A(\router/ram_read_enable_reg ));
   CLKBUFX2TS FE_OFC1283_router_fft_write_done (.Y(FE_OFN1283_router_fft_write_done), 
	.A(\router/fft_write_done ));
   CLKBUFX2TS FE_OFC1282_router_fft_get_req_reg (.Y(FE_OFN1282_router_fft_get_req_reg), 
	.A(\router/fft_get_req_reg ));
   CLKBUFX2TS FE_OFC1281_router_addr_calc_iir_write_calc_count_5_ (.Y(FE_OFN1281_router_addr_calc_iir_write_calc_count_5_), 
	.A(\router/addr_calc/iir_write_calc/count[5] ));
   CLKBUFX2TS FE_OFC1280_router_addr_calc_iir_write_calc_count_9_ (.Y(FE_OFN1280_router_addr_calc_iir_write_calc_count_9_), 
	.A(\router/addr_calc/iir_write_calc/count[9] ));
   CLKBUFX2TS FE_OFC1279_n7328 (.Y(FE_OFN1279_n7328), 
	.A(n7328));
   CLKBUFX2TS FE_OFC1278_n7333 (.Y(FE_OFN1278_n7333), 
	.A(n7333));
   CLKBUFX2TS FE_OFC1277_n7308 (.Y(FE_OFN1277_n7308), 
	.A(n7308));
   CLKBUFX2TS FE_OFC1276_router_addr_calc_fir_read_calc_count_5_ (.Y(FE_OFN1276_router_addr_calc_fir_read_calc_count_5_), 
	.A(FE_OFN1824_router_addr_calc_fir_read_calc_count_5_));
   CLKBUFX2TS FE_OFC1275_n7353 (.Y(FE_OFN1275_n7353), 
	.A(n7353));
   CLKBUFX2TS FE_OFC1274_n7358 (.Y(FE_OFN1274_n7358), 
	.A(n7358));
   CLKBUFX2TS FE_OFC1273_router_addr_calc_fft_read_calc_count_5_ (.Y(FE_OFN1273_router_addr_calc_fft_read_calc_count_5_), 
	.A(\router/addr_calc/fft_read_calc/count[5] ));
   CLKBUFX2TS FE_OFC1272_router_addr_calc_fir_write_calc_count_5_ (.Y(FE_OFN1272_router_addr_calc_fir_write_calc_count_5_), 
	.A(\router/addr_calc/fir_write_calc/count[5] ));
   CLKBUFX2TS FE_OFC1271_router_addr_calc_fir_read_calc_count_15_ (.Y(FE_OFN1271_router_addr_calc_fir_read_calc_count_15_), 
	.A(\router/addr_calc/fir_read_calc/count[15] ));
   CLKBUFX2TS FE_OFC1270_router_addr_calc_fft_write_calc_count_15_ (.Y(FE_OFN1270_router_addr_calc_fft_write_calc_count_15_), 
	.A(\router/addr_calc/fft_write_calc/count[15] ));
   CLKBUFX2TS FE_OFC1269_router_addr_calc_fir_read_calc_count_9_ (.Y(FE_OFN1269_router_addr_calc_fir_read_calc_count_9_), 
	.A(\router/addr_calc/fir_read_calc/count[9] ));
   CLKBUFX2TS FE_OFC1268_router_addr_calc_fft_write_calc_count_9_ (.Y(FE_OFN1268_router_addr_calc_fft_write_calc_count_9_), 
	.A(\router/addr_calc/fft_write_calc/count[9] ));
   CLKBUFX2TS FE_OFC1267_router_addr_calc_fft_read_calc_count_9_ (.Y(FE_OFN1267_router_addr_calc_fft_read_calc_count_9_), 
	.A(\router/addr_calc/fft_read_calc/count[9] ));
   CLKBUFX2TS FE_OFC1266_router_addr_calc_fir_write_calc_count_9_ (.Y(FE_OFN1266_router_addr_calc_fir_write_calc_count_9_), 
	.A(\router/addr_calc/fir_write_calc/count[9] ));
   CLKBUFX2TS FE_OFC1265_n7303 (.Y(FE_OFN1265_n7303), 
	.A(n7303));
   CLKBUFX2TS FE_OFC1264_router_addr_calc_fir_write_calc_count_16_ (.Y(FE_OFN1264_router_addr_calc_fir_write_calc_count_16_), 
	.A(\router/addr_calc/fir_write_calc/count[16] ));
   CLKBUFX2TS FE_OFC1263_router_addr_calc_fft_read_calc_count_16_ (.Y(FE_OFN1263_router_addr_calc_fft_read_calc_count_16_), 
	.A(\router/addr_calc/fft_read_calc/count[16] ));
   CLKBUFX2TS FE_OFC1262_n7298 (.Y(FE_OFN1262_n7298), 
	.A(n7298));
   CLKBUFX2TS FE_OFC1261_router_addr_calc_fir_write_calc_count_19_ (.Y(FE_OFN1261_router_addr_calc_fir_write_calc_count_19_), 
	.A(\router/addr_calc/fir_write_calc/count[19] ));
   CLKBUFX2TS FE_OFC1260_router_addr_calc_fir_read_calc_count_19_ (.Y(FE_OFN1260_router_addr_calc_fir_read_calc_count_19_), 
	.A(\router/addr_calc/fir_read_calc/count[19] ));
   CLKBUFX2TS FE_OFC1259_router_addr_calc_fft_write_calc_count_19_ (.Y(FE_OFN1259_router_addr_calc_fft_write_calc_count_19_), 
	.A(\router/addr_calc/fft_write_calc/count[19] ));
   CLKBUFX2TS FE_OFC1258_router_addr_calc_fft_read_calc_count_19_ (.Y(FE_OFN1258_router_addr_calc_fft_read_calc_count_19_), 
	.A(\router/addr_calc/fft_read_calc/count[19] ));
   CLKBUFX2TS FE_OFC1257_n7165 (.Y(FE_OFN1257_n7165), 
	.A(n7165));
   CLKBUFX2TS FE_OFC1256_n7288 (.Y(FE_OFN1256_n7288), 
	.A(n7288));
   CLKBUFX2TS FE_OFC1255_n7402 (.Y(FE_OFN1255_n7402), 
	.A(n7402));
   CLKBUFX2TS FE_OFC1254_n7159 (.Y(FE_OFN1254_n7159), 
	.A(n7159));
   CLKBUFX2TS FE_OFC1253_n7283 (.Y(FE_OFN1253_n7283), 
	.A(n7283));
   CLKBUFX2TS FE_OFC1252_n7397 (.Y(FE_OFN1252_n7397), 
	.A(n7397));
   CLKBUFX2TS FE_OFC1251_n7153 (.Y(FE_OFN1251_n7153), 
	.A(n7153));
   CLKBUFX2TS FE_OFC1250_n7278 (.Y(FE_OFN1250_n7278), 
	.A(n7278));
   CLKBUFX2TS FE_OFC1249_n7392 (.Y(FE_OFN1249_n7392), 
	.A(n7392));
   CLKBUFX2TS FE_OFC1248_router_addr_calc_fir_write_calc_count_23_ (.Y(FE_OFN1248_router_addr_calc_fir_write_calc_count_23_), 
	.A(\router/addr_calc/fir_write_calc/count[23] ));
   CLKBUFX2TS FE_OFC1247_router_addr_calc_fir_read_calc_count_23_ (.Y(FE_OFN1247_router_addr_calc_fir_read_calc_count_23_), 
	.A(\router/addr_calc/fir_read_calc/count[23] ));
   CLKBUFX2TS FE_OFC1246_router_addr_calc_fft_write_calc_count_23_ (.Y(FE_OFN1246_router_addr_calc_fft_write_calc_count_23_), 
	.A(\router/addr_calc/fft_write_calc/count[23] ));
   CLKBUFX2TS FE_OFC1245_router_addr_calc_fft_read_calc_count_23_ (.Y(FE_OFN1245_router_addr_calc_fft_read_calc_count_23_), 
	.A(\router/addr_calc/fft_read_calc/count[23] ));
   CLKBUFX2TS FE_OFC1244_router_addr_calc_iir_write_calc_count_23_ (.Y(FE_OFN1244_router_addr_calc_iir_write_calc_count_23_), 
	.A(\router/addr_calc/iir_write_calc/count[23] ));
   CLKBUFX2TS FE_OFC1243_n7273 (.Y(FE_OFN1243_n7273), 
	.A(n7273));
   CLKBUFX2TS FE_OFC1242_n7268 (.Y(FE_OFN1242_n7268), 
	.A(n7268));
   CLKBUFX2TS FE_OFC1241_n7264 (.Y(FE_OFN1241_n7264), 
	.A(n7264));
   CLKBUFX2TS FE_OFC1240_router_addr_calc_fir_write_calc_count_27_ (.Y(FE_OFN1240_router_addr_calc_fir_write_calc_count_27_), 
	.A(\router/addr_calc/fir_write_calc/count[27] ));
   CLKBUFX2TS FE_OFC1239_router_addr_calc_fir_read_calc_count_27_ (.Y(FE_OFN1239_router_addr_calc_fir_read_calc_count_27_), 
	.A(\router/addr_calc/fir_read_calc/count[27] ));
   CLKBUFX2TS FE_OFC1238_router_addr_calc_fft_write_calc_count_27_ (.Y(FE_OFN1238_router_addr_calc_fft_write_calc_count_27_), 
	.A(\router/addr_calc/fft_write_calc/count[27] ));
   CLKBUFX2TS FE_OFC1237_router_addr_calc_fft_read_calc_count_27_ (.Y(FE_OFN1237_router_addr_calc_fft_read_calc_count_27_), 
	.A(\router/addr_calc/fft_read_calc/count[27] ));
   CLKBUFX2TS FE_OFC1236_n7259 (.Y(FE_OFN1236_n7259), 
	.A(n7259));
   CLKBUFX2TS FE_OFC1235_n7254 (.Y(FE_OFN1235_n7254), 
	.A(n7254));
   CLKBUFX2TS FE_OFC1234_n7492 (.Y(FE_OFN1234_n7492), 
	.A(n7492));
   CLKBUFX2TS FE_OFC1233_router_addr_calc_fft_write_calc_count_29_ (.Y(FE_OFN1233_router_addr_calc_fft_write_calc_count_29_), 
	.A(\router/addr_calc/fft_write_calc/count[29] ));
   CLKBUFX2TS FE_OFC1232_n7368 (.Y(FE_OFN1232_n7368), 
	.A(n7368));
   CLKBUFX2TS FE_OFC1231_router_addr_calc_fir_write_calc_count_30_ (.Y(FE_OFN1231_router_addr_calc_fir_write_calc_count_30_), 
	.A(\router/addr_calc/fir_write_calc/count[30] ));
   CLKBUFX2TS FE_OFC1230_router_addr_calc_fir_read_calc_count_30_ (.Y(FE_OFN1230_router_addr_calc_fir_read_calc_count_30_), 
	.A(\router/addr_calc/fir_read_calc/count[30] ));
   CLKBUFX2TS FE_OFC1229_router_addr_calc_fft_read_calc_count_30_ (.Y(FE_OFN1229_router_addr_calc_fft_read_calc_count_30_), 
	.A(\router/addr_calc/fft_read_calc/count[30] ));
   CLKBUFX2TS FE_OFC1228_router_addr_calc_fft_write_calc_count_31_ (.Y(FE_OFN1228_router_addr_calc_fft_write_calc_count_31_), 
	.A(\router/addr_calc/fft_write_calc/count[31] ));
   CLKBUFX2TS FE_OFC1227_n8063 (.Y(FE_OFN1227_n8063), 
	.A(FE_OFN1226_n8063));
   CLKBUFX2TS FE_OFC1226_n8063 (.Y(FE_OFN1226_n8063), 
	.A(FE_OFN1225_n8063));
   CLKBUFX2TS FE_OFC1225_n8063 (.Y(FE_OFN1225_n8063), 
	.A(FE_OFN1223_n8063));
   CLKBUFX2TS FE_OFC1224_n8063 (.Y(FE_OFN1224_n8063), 
	.A(n8063));
   CLKBUFX2TS FE_OFC1223_n8063 (.Y(FE_OFN1223_n8063), 
	.A(n8063));
   CLKBUFX2TS FE_OFC1222_n8064 (.Y(FE_OFN1222_n8064), 
	.A(FE_OFN1221_n8064));
   CLKBUFX2TS FE_OFC1221_n8064 (.Y(FE_OFN1221_n8064), 
	.A(FE_OFN1219_n8064));
   CLKBUFX2TS FE_OFC1220_n8064 (.Y(FE_OFN1220_n8064), 
	.A(FE_OFN1219_n8064));
   CLKBUFX2TS FE_OFC1219_n8064 (.Y(FE_OFN1219_n8064), 
	.A(FE_OFN1218_n8064));
   CLKBUFX2TS FE_OFC1218_n8064 (.Y(FE_OFN1218_n8064), 
	.A(n8064));
   CLKBUFX2TS FE_OFC1217_n3478 (.Y(FE_OFN1217_n3478), 
	.A(n3478));
   CLKBUFX2TS FE_OFC1216_n8061 (.Y(FE_OFN1216_n8061), 
	.A(FE_OFN1215_n8061));
   CLKBUFX2TS FE_OFC1215_n8061 (.Y(FE_OFN1215_n8061), 
	.A(FE_OFN1214_n8061));
   CLKBUFX2TS FE_OFC1214_n8061 (.Y(FE_OFN1214_n8061), 
	.A(FE_OFN1212_n8061));
   CLKBUFX2TS FE_OFC1213_n8061 (.Y(FE_OFN1213_n8061), 
	.A(FE_OFN1212_n8061));
   CLKBUFX2TS FE_OFC1212_n8061 (.Y(FE_OFN1212_n8061), 
	.A(n8061));
   CLKBUFX2TS FE_OFC1211_n8062 (.Y(FE_OFN1211_n8062), 
	.A(FE_OFN1209_n8062));
   CLKBUFX2TS FE_OFC1210_n8062 (.Y(FE_OFN1210_n8062), 
	.A(FE_OFN1209_n8062));
   CLKBUFX2TS FE_OFC1209_n8062 (.Y(FE_OFN1209_n8062), 
	.A(FE_OFN1208_n8062));
   CLKBUFX2TS FE_OFC1208_n8062 (.Y(FE_OFN1208_n8062), 
	.A(n8062));
   CLKBUFX2TS FE_OFC1207_router_addr_calc_iir_write_calc_counter_N212 (.Y(FE_OFN1207_router_addr_calc_iir_write_calc_counter_N212), 
	.A(FE_OFN1206_router_addr_calc_iir_write_calc_counter_N212));
   CLKBUFX2TS FE_OFC1206_router_addr_calc_iir_write_calc_counter_N212 (.Y(FE_OFN1206_router_addr_calc_iir_write_calc_counter_N212), 
	.A(FE_OFN1204_router_addr_calc_iir_write_calc_counter_N212));
   CLKBUFX2TS FE_OFC1205_router_addr_calc_iir_write_calc_counter_N212 (.Y(FE_OFN1205_router_addr_calc_iir_write_calc_counter_N212), 
	.A(FE_OFN1203_router_addr_calc_iir_write_calc_counter_N212));
   CLKBUFX2TS FE_OFC1204_router_addr_calc_iir_write_calc_counter_N212 (.Y(FE_OFN1204_router_addr_calc_iir_write_calc_counter_N212), 
	.A(FE_OFN1203_router_addr_calc_iir_write_calc_counter_N212));
   CLKBUFX2TS FE_OFC1203_router_addr_calc_iir_write_calc_counter_N212 (.Y(FE_OFN1203_router_addr_calc_iir_write_calc_counter_N212), 
	.A(FE_OFN1202_router_addr_calc_iir_write_calc_counter_N212));
   CLKBUFX2TS FE_OFC1202_router_addr_calc_iir_write_calc_counter_N212 (.Y(FE_OFN1202_router_addr_calc_iir_write_calc_counter_N212), 
	.A(FE_OFN1201_router_addr_calc_iir_write_calc_counter_N212));
   CLKBUFX2TS FE_OFC1201_router_addr_calc_iir_write_calc_counter_N212 (.Y(FE_OFN1201_router_addr_calc_iir_write_calc_counter_N212), 
	.A(FE_OFN1200_router_addr_calc_iir_write_calc_counter_N212));
   CLKBUFX2TS FE_OFC1200_router_addr_calc_iir_write_calc_counter_N212 (.Y(FE_OFN1200_router_addr_calc_iir_write_calc_counter_N212), 
	.A(FE_OFN1199_router_addr_calc_iir_write_calc_counter_N212));
   CLKBUFX2TS FE_OFC1199_router_addr_calc_iir_write_calc_counter_N212 (.Y(FE_OFN1199_router_addr_calc_iir_write_calc_counter_N212), 
	.A(\router/addr_calc/iir_write_calc/counter/N212 ));
   CLKBUFX2TS FE_OFC1198_n7023 (.Y(FE_OFN1198_n7023), 
	.A(FE_OFN1197_n7023));
   CLKBUFX2TS FE_OFC1197_n7023 (.Y(FE_OFN1197_n7023), 
	.A(FE_OFN1196_n7023));
   CLKBUFX2TS FE_OFC1196_n7023 (.Y(FE_OFN1196_n7023), 
	.A(FE_OFN1195_n7023));
   CLKBUFX2TS FE_OFC1195_n7023 (.Y(FE_OFN1195_n7023), 
	.A(FE_OFN1194_n7023));
   CLKBUFX2TS FE_OFC1194_n7023 (.Y(FE_OFN1194_n7023), 
	.A(FE_OFN1193_n7023));
   CLKBUFX2TS FE_OFC1193_n7023 (.Y(FE_OFN1193_n7023), 
	.A(n7023));
   CLKBUFX2TS FE_OFC1192_n7022 (.Y(FE_OFN1192_n7022), 
	.A(FE_OFN1190_n7022));
   CLKBUFX2TS FE_OFC1191_n7022 (.Y(FE_OFN1191_n7022), 
	.A(n7022));
   CLKBUFX2TS FE_OFC1190_n7022 (.Y(FE_OFN1190_n7022), 
	.A(n7022));
   CLKBUFX2TS FE_OFC1189_n7020 (.Y(FE_OFN1189_n7020), 
	.A(FE_OFN1186_n7020));
   CLKBUFX2TS FE_OFC1188_n7020 (.Y(FE_OFN1188_n7020), 
	.A(FE_OFN1187_n7020));
   CLKBUFX2TS FE_OFC1187_n7020 (.Y(FE_OFN1187_n7020), 
	.A(FE_OFN1184_n7020));
   CLKBUFX2TS FE_OFC1186_n7020 (.Y(FE_OFN1186_n7020), 
	.A(FE_OFN1185_n7020));
   CLKBUFX2TS FE_OFC1185_n7020 (.Y(FE_OFN1185_n7020), 
	.A(FE_OFN1182_n7020));
   CLKBUFX2TS FE_OFC1184_n7020 (.Y(FE_OFN1184_n7020), 
	.A(FE_OFN1183_n7020));
   CLKBUFX2TS FE_OFC1183_n7020 (.Y(FE_OFN1183_n7020), 
	.A(FE_OFN1181_n7020));
   CLKBUFX2TS FE_OFC1182_n7020 (.Y(FE_OFN1182_n7020), 
	.A(FE_OFN1180_n7020));
   CLKBUFX2TS FE_OFC1181_n7020 (.Y(FE_OFN1181_n7020), 
	.A(FE_OFN1180_n7020));
   CLKBUFX2TS FE_OFC1180_n7020 (.Y(FE_OFN1180_n7020), 
	.A(FE_OFN1179_n7020));
   CLKBUFX2TS FE_OFC1179_n7020 (.Y(FE_OFN1179_n7020), 
	.A(n7020));
   CLKBUFX2TS FE_OFC1178_n7021 (.Y(FE_OFN1178_n7021), 
	.A(FE_OFN1176_n7021));
   CLKBUFX2TS FE_OFC1177_n7021 (.Y(FE_OFN1177_n7021), 
	.A(FE_OFN1175_n7021));
   CLKBUFX2TS FE_OFC1176_n7021 (.Y(FE_OFN1176_n7021), 
	.A(FE_OFN1174_n7021));
   CLKBUFX2TS FE_OFC1175_n7021 (.Y(FE_OFN1175_n7021), 
	.A(FE_OFN1174_n7021));
   CLKBUFX2TS FE_OFC1174_n7021 (.Y(FE_OFN1174_n7021), 
	.A(FE_OFN1172_n7021));
   CLKBUFX2TS FE_OFC1173_n7021 (.Y(FE_OFN1173_n7021), 
	.A(FE_OFN1172_n7021));
   CLKBUFX2TS FE_OFC1172_n7021 (.Y(FE_OFN1172_n7021), 
	.A(FE_OFN1171_n7021));
   CLKBUFX2TS FE_OFC1171_n7021 (.Y(FE_OFN1171_n7021), 
	.A(FE_OFN1168_n7021));
   CLKBUFX2TS FE_OFC1170_n7021 (.Y(FE_OFN1170_n7021), 
	.A(FE_OFN1169_n7021));
   CLKBUFX2TS FE_OFC1169_n7021 (.Y(FE_OFN1169_n7021), 
	.A(n7021));
   CLKBUFX2TS FE_OFC1168_n7021 (.Y(FE_OFN1168_n7021), 
	.A(n7021));
   CLKBUFX2TS FE_OFC1167_n7019 (.Y(FE_OFN1167_n7019), 
	.A(FE_OFN1164_n7019));
   CLKBUFX2TS FE_OFC1166_n7019 (.Y(FE_OFN1166_n7019), 
	.A(FE_OFN1163_n7019));
   CLKBUFX2TS FE_OFC1165_n7019 (.Y(FE_OFN1165_n7019), 
	.A(FE_OFN1163_n7019));
   CLKBUFX2TS FE_OFC1164_n7019 (.Y(FE_OFN1164_n7019), 
	.A(FE_OFN1162_n7019));
   CLKBUFX2TS FE_OFC1163_n7019 (.Y(FE_OFN1163_n7019), 
	.A(FE_OFN1160_n7019));
   CLKBUFX2TS FE_OFC1162_n7019 (.Y(FE_OFN1162_n7019), 
	.A(FE_OFN1161_n7019));
   CLKBUFX2TS FE_OFC1161_n7019 (.Y(FE_OFN1161_n7019), 
	.A(FE_OFN1159_n7019));
   CLKBUFX2TS FE_OFC1160_n7019 (.Y(FE_OFN1160_n7019), 
	.A(FE_OFN1159_n7019));
   CLKBUFX2TS FE_OFC1159_n7019 (.Y(FE_OFN1159_n7019), 
	.A(FE_OFN1158_n7019));
   CLKBUFX2TS FE_OFC1158_n7019 (.Y(FE_OFN1158_n7019), 
	.A(n7019));
   CLKBUFX2TS FE_OFC1157_n1609 (.Y(FE_OFN1157_n1609), 
	.A(FE_OFN1155_n1609));
   CLKBUFX2TS FE_OFC1156_n1609 (.Y(FE_OFN1156_n1609), 
	.A(FE_OFN1154_n1609));
   CLKBUFX2TS FE_OFC1155_n1609 (.Y(FE_OFN1155_n1609), 
	.A(FE_OFN1153_n1609));
   CLKBUFX2TS FE_OFC1154_n1609 (.Y(FE_OFN1154_n1609), 
	.A(FE_OFN1152_n1609));
   CLKBUFX2TS FE_OFC1153_n1609 (.Y(FE_OFN1153_n1609), 
	.A(FE_OFN1152_n1609));
   CLKBUFX2TS FE_OFC1152_n1609 (.Y(FE_OFN1152_n1609), 
	.A(FE_OFN1151_n1609));
   CLKBUFX2TS FE_OFC1151_n1609 (.Y(FE_OFN1151_n1609), 
	.A(FE_OFN1149_n1609));
   CLKBUFX2TS FE_OFC1150_n1609 (.Y(FE_OFN1150_n1609), 
	.A(FE_OFN1149_n1609));
   CLKBUFX2TS FE_OFC1149_n1609 (.Y(FE_OFN1149_n1609), 
	.A(FE_OFN1148_n1609));
   CLKBUFX2TS FE_OFC1148_n1609 (.Y(FE_OFN1148_n1609), 
	.A(n1609));
   CLKBUFX2TS FE_OFC1147_n585 (.Y(FE_OFN1147_n585), 
	.A(FE_OFN1146_n585));
   CLKBUFX2TS FE_OFC1146_n585 (.Y(FE_OFN1146_n585), 
	.A(FE_OFN1145_n585));
   CLKBUFX2TS FE_OFC1145_n585 (.Y(FE_OFN1145_n585), 
	.A(FE_OFN1142_n585));
   CLKBUFX2TS FE_OFC1144_n585 (.Y(FE_OFN1144_n585), 
	.A(FE_OFN1140_n585));
   CLKBUFX2TS FE_OFC1143_n585 (.Y(FE_OFN1143_n585), 
	.A(FE_OFN1141_n585));
   CLKBUFX2TS FE_OFC1142_n585 (.Y(FE_OFN1142_n585), 
	.A(FE_OFN1140_n585));
   CLKBUFX2TS FE_OFC1141_n585 (.Y(FE_OFN1141_n585), 
	.A(FE_OFN1138_n585));
   CLKBUFX2TS FE_OFC1140_n585 (.Y(FE_OFN1140_n585), 
	.A(FE_OFN1139_n585));
   CLKBUFX2TS FE_OFC1139_n585 (.Y(FE_OFN1139_n585), 
	.A(FE_OFN1138_n585));
   CLKBUFX2TS FE_OFC1138_n585 (.Y(FE_OFN1138_n585), 
	.A(n585));
   CLKBUFX2TS FE_OFC1137_n2505 (.Y(FE_OFN1137_n2505), 
	.A(FE_OFN1136_n2505));
   CLKBUFX2TS FE_OFC1136_n2505 (.Y(FE_OFN1136_n2505), 
	.A(FE_OFN1134_n2505));
   CLKBUFX2TS FE_OFC1135_n2505 (.Y(FE_OFN1135_n2505), 
	.A(FE_OFN1133_n2505));
   CLKBUFX2TS FE_OFC1134_n2505 (.Y(FE_OFN1134_n2505), 
	.A(FE_OFN1133_n2505));
   CLKBUFX2TS FE_OFC1133_n2505 (.Y(FE_OFN1133_n2505), 
	.A(n2505));
   CLKBUFX2TS FE_OFC1132_n2441 (.Y(FE_OFN1132_n2441), 
	.A(FE_OFN1130_n2441));
   CLKBUFX2TS FE_OFC1131_n2441 (.Y(FE_OFN1131_n2441), 
	.A(FE_OFN1130_n2441));
   CLKBUFX2TS FE_OFC1130_n2441 (.Y(FE_OFN1130_n2441), 
	.A(FE_OFN1129_n2441));
   CLKBUFX2TS FE_OFC1129_n2441 (.Y(FE_OFN1129_n2441), 
	.A(n2441));
   CLKBUFX2TS FE_OFC1128_n2377 (.Y(FE_OFN1128_n2377), 
	.A(FE_OFN1126_n2377));
   CLKBUFX2TS FE_OFC1127_n2377 (.Y(FE_OFN1127_n2377), 
	.A(FE_OFN1126_n2377));
   CLKBUFX2TS FE_OFC1126_n2377 (.Y(FE_OFN1126_n2377), 
	.A(FE_OFN1125_n2377));
   CLKBUFX2TS FE_OFC1125_n2377 (.Y(FE_OFN1125_n2377), 
	.A(FE_OFN1124_n2377));
   CLKBUFX2TS FE_OFC1124_n2377 (.Y(FE_OFN1124_n2377), 
	.A(n2377));
   CLKBUFX2TS FE_OFC1123_n2313 (.Y(FE_OFN1123_n2313), 
	.A(FE_OFN1122_n2313));
   CLKBUFX2TS FE_OFC1122_n2313 (.Y(FE_OFN1122_n2313), 
	.A(FE_OFN1121_n2313));
   CLKBUFX2TS FE_OFC1121_n2313 (.Y(FE_OFN1121_n2313), 
	.A(FE_OFN1120_n2313));
   CLKBUFX2TS FE_OFC1120_n2313 (.Y(FE_OFN1120_n2313), 
	.A(n2313));
   CLKBUFX2TS FE_OFC1119_n2249 (.Y(FE_OFN1119_n2249), 
	.A(FE_OFN1117_n2249));
   CLKBUFX2TS FE_OFC1118_n2249 (.Y(FE_OFN1118_n2249), 
	.A(FE_OFN1117_n2249));
   CLKBUFX2TS FE_OFC1117_n2249 (.Y(FE_OFN1117_n2249), 
	.A(FE_OFN1116_n2249));
   CLKBUFX2TS FE_OFC1116_n2249 (.Y(FE_OFN1116_n2249), 
	.A(FE_OFN1115_n2249));
   CLKBUFX2TS FE_OFC1115_n2249 (.Y(FE_OFN1115_n2249), 
	.A(n2249));
   CLKBUFX2TS FE_OFC1114_n2185 (.Y(FE_OFN1114_n2185), 
	.A(FE_OFN1112_n2185));
   CLKBUFX2TS FE_OFC1113_n2185 (.Y(FE_OFN1113_n2185), 
	.A(FE_OFN1111_n2185));
   CLKBUFX2TS FE_OFC1112_n2185 (.Y(FE_OFN1112_n2185), 
	.A(n2185));
   CLKBUFX2TS FE_OFC1111_n2185 (.Y(FE_OFN1111_n2185), 
	.A(n2185));
   CLKBUFX2TS FE_OFC1110_n2121 (.Y(FE_OFN1110_n2121), 
	.A(FE_OFN1107_n2121));
   CLKBUFX2TS FE_OFC1109_n2121 (.Y(FE_OFN1109_n2121), 
	.A(FE_OFN1106_n2121));
   CLKBUFX2TS FE_OFC1108_n2121 (.Y(FE_OFN1108_n2121), 
	.A(FE_OFN1107_n2121));
   CLKBUFX2TS FE_OFC1107_n2121 (.Y(FE_OFN1107_n2121), 
	.A(FE_OFN1106_n2121));
   CLKBUFX2TS FE_OFC1106_n2121 (.Y(FE_OFN1106_n2121), 
	.A(n2121));
   CLKBUFX2TS FE_OFC1105_n2057 (.Y(FE_OFN1105_n2057), 
	.A(FE_OFN1104_n2057));
   CLKBUFX2TS FE_OFC1104_n2057 (.Y(FE_OFN1104_n2057), 
	.A(FE_OFN1103_n2057));
   CLKBUFX2TS FE_OFC1103_n2057 (.Y(FE_OFN1103_n2057), 
	.A(FE_OFN1102_n2057));
   CLKBUFX2TS FE_OFC1102_n2057 (.Y(FE_OFN1102_n2057), 
	.A(n2057));
   CLKBUFX2TS FE_OFC1101_n1993 (.Y(FE_OFN1101_n1993), 
	.A(FE_OFN1100_n1993));
   CLKBUFX2TS FE_OFC1100_n1993 (.Y(FE_OFN1100_n1993), 
	.A(FE_OFN1098_n1993));
   CLKBUFX2TS FE_OFC1099_n1993 (.Y(FE_OFN1099_n1993), 
	.A(FE_OFN1097_n1993));
   CLKBUFX2TS FE_OFC1098_n1993 (.Y(FE_OFN1098_n1993), 
	.A(FE_OFN1097_n1993));
   CLKBUFX2TS FE_OFC1097_n1993 (.Y(FE_OFN1097_n1993), 
	.A(n1993));
   CLKBUFX2TS FE_OFC1096_n1929 (.Y(FE_OFN1096_n1929), 
	.A(FE_OFN1095_n1929));
   CLKBUFX2TS FE_OFC1095_n1929 (.Y(FE_OFN1095_n1929), 
	.A(FE_OFN1094_n1929));
   CLKBUFX2TS FE_OFC1094_n1929 (.Y(FE_OFN1094_n1929), 
	.A(FE_OFN1093_n1929));
   CLKBUFX2TS FE_OFC1093_n1929 (.Y(FE_OFN1093_n1929), 
	.A(n1929));
   CLKBUFX2TS FE_OFC1092_n1865 (.Y(FE_OFN1092_n1865), 
	.A(FE_OFN1091_n1865));
   CLKBUFX2TS FE_OFC1091_n1865 (.Y(FE_OFN1091_n1865), 
	.A(FE_OFN1090_n1865));
   CLKBUFX2TS FE_OFC1090_n1865 (.Y(FE_OFN1090_n1865), 
	.A(FE_OFN1089_n1865));
   CLKBUFX2TS FE_OFC1089_n1865 (.Y(FE_OFN1089_n1865), 
	.A(n1865));
   CLKBUFX2TS FE_OFC1088_n1801 (.Y(FE_OFN1088_n1801), 
	.A(FE_OFN1087_n1801));
   CLKBUFX2TS FE_OFC1087_n1801 (.Y(FE_OFN1087_n1801), 
	.A(FE_OFN1086_n1801));
   CLKBUFX2TS FE_OFC1086_n1801 (.Y(FE_OFN1086_n1801), 
	.A(FE_OFN1085_n1801));
   CLKBUFX2TS FE_OFC1085_n1801 (.Y(FE_OFN1085_n1801), 
	.A(n1801));
   CLKBUFX2TS FE_OFC1084_n1737 (.Y(FE_OFN1084_n1737), 
	.A(FE_OFN1081_n1737));
   CLKBUFX2TS FE_OFC1083_n1737 (.Y(FE_OFN1083_n1737), 
	.A(FE_OFN1081_n1737));
   CLKBUFX2TS FE_OFC1082_n1737 (.Y(FE_OFN1082_n1737), 
	.A(n1737));
   CLKBUFX2TS FE_OFC1081_n1737 (.Y(FE_OFN1081_n1737), 
	.A(n1737));
   CLKBUFX2TS FE_OFC1080_n1673 (.Y(FE_OFN1080_n1673), 
	.A(FE_OFN1078_n1673));
   CLKBUFX2TS FE_OFC1079_n1673 (.Y(FE_OFN1079_n1673), 
	.A(FE_OFN1077_n1673));
   CLKBUFX2TS FE_OFC1078_n1673 (.Y(FE_OFN1078_n1673), 
	.A(FE_OFN1077_n1673));
   CLKBUFX2TS FE_OFC1077_n1673 (.Y(FE_OFN1077_n1673), 
	.A(n1673));
   CLKBUFX2TS FE_OFC1076_n1481 (.Y(FE_OFN1076_n1481), 
	.A(FE_OFN1075_n1481));
   CLKBUFX2TS FE_OFC1075_n1481 (.Y(FE_OFN1075_n1481), 
	.A(FE_OFN1074_n1481));
   CLKBUFX2TS FE_OFC1074_n1481 (.Y(FE_OFN1074_n1481), 
	.A(FE_OFN1073_n1481));
   CLKBUFX2TS FE_OFC1073_n1481 (.Y(FE_OFN1073_n1481), 
	.A(n1481));
   CLKBUFX2TS FE_OFC1072_n1417 (.Y(FE_OFN1072_n1417), 
	.A(FE_OFN1071_n1417));
   CLKBUFX2TS FE_OFC1071_n1417 (.Y(FE_OFN1071_n1417), 
	.A(FE_OFN1070_n1417));
   CLKBUFX2TS FE_OFC1070_n1417 (.Y(FE_OFN1070_n1417), 
	.A(FE_OFN1069_n1417));
   CLKBUFX2TS FE_OFC1069_n1417 (.Y(FE_OFN1069_n1417), 
	.A(n1417));
   CLKBUFX2TS FE_OFC1068_n1353 (.Y(FE_OFN1068_n1353), 
	.A(FE_OFN1067_n1353));
   CLKBUFX2TS FE_OFC1067_n1353 (.Y(FE_OFN1067_n1353), 
	.A(FE_OFN1066_n1353));
   CLKBUFX2TS FE_OFC1066_n1353 (.Y(FE_OFN1066_n1353), 
	.A(n1353));
   CLKBUFX2TS FE_OFC1065_n1353 (.Y(FE_OFN1065_n1353), 
	.A(n1353));
   CLKBUFX2TS FE_OFC1064_n1289 (.Y(FE_OFN1064_n1289), 
	.A(FE_OFN1063_n1289));
   CLKBUFX2TS FE_OFC1063_n1289 (.Y(FE_OFN1063_n1289), 
	.A(FE_OFN1062_n1289));
   CLKBUFX2TS FE_OFC1062_n1289 (.Y(FE_OFN1062_n1289), 
	.A(FE_OFN1061_n1289));
   CLKBUFX2TS FE_OFC1061_n1289 (.Y(FE_OFN1061_n1289), 
	.A(n1289));
   CLKBUFX2TS FE_OFC1060_n1225 (.Y(FE_OFN1060_n1225), 
	.A(FE_OFN1059_n1225));
   CLKBUFX2TS FE_OFC1059_n1225 (.Y(FE_OFN1059_n1225), 
	.A(FE_OFN1058_n1225));
   CLKBUFX2TS FE_OFC1058_n1225 (.Y(FE_OFN1058_n1225), 
	.A(FE_OFN1057_n1225));
   CLKBUFX2TS FE_OFC1057_n1225 (.Y(FE_OFN1057_n1225), 
	.A(FE_OFN1056_n1225));
   CLKBUFX2TS FE_OFC1056_n1225 (.Y(FE_OFN1056_n1225), 
	.A(n1225));
   CLKBUFX2TS FE_OFC1055_n1161 (.Y(FE_OFN1055_n1161), 
	.A(FE_OFN1054_n1161));
   CLKBUFX2TS FE_OFC1054_n1161 (.Y(FE_OFN1054_n1161), 
	.A(FE_OFN1053_n1161));
   CLKBUFX2TS FE_OFC1053_n1161 (.Y(FE_OFN1053_n1161), 
	.A(FE_OFN1052_n1161));
   CLKBUFX2TS FE_OFC1052_n1161 (.Y(FE_OFN1052_n1161), 
	.A(n1161));
   CLKBUFX2TS FE_OFC1051_n1097 (.Y(FE_OFN1051_n1097), 
	.A(FE_OFN1050_n1097));
   CLKBUFX2TS FE_OFC1050_n1097 (.Y(FE_OFN1050_n1097), 
	.A(FE_OFN1049_n1097));
   CLKBUFX2TS FE_OFC1049_n1097 (.Y(FE_OFN1049_n1097), 
	.A(FE_OFN1048_n1097));
   CLKBUFX2TS FE_OFC1048_n1097 (.Y(FE_OFN1048_n1097), 
	.A(n1097));
   CLKBUFX2TS FE_OFC1047_n1033 (.Y(FE_OFN1047_n1033), 
	.A(FE_OFN1046_n1033));
   CLKBUFX2TS FE_OFC1046_n1033 (.Y(FE_OFN1046_n1033), 
	.A(FE_OFN1044_n1033));
   CLKBUFX2TS FE_OFC1045_n1033 (.Y(FE_OFN1045_n1033), 
	.A(FE_OFN1044_n1033));
   CLKBUFX2TS FE_OFC1044_n1033 (.Y(FE_OFN1044_n1033), 
	.A(FE_OFN1043_n1033));
   CLKBUFX2TS FE_OFC1043_n1033 (.Y(FE_OFN1043_n1033), 
	.A(n1033));
   CLKBUFX2TS FE_OFC1042_n969 (.Y(FE_OFN1042_n969), 
	.A(FE_OFN1041_n969));
   CLKBUFX2TS FE_OFC1041_n969 (.Y(FE_OFN1041_n969), 
	.A(FE_OFN1040_n969));
   CLKBUFX2TS FE_OFC1040_n969 (.Y(FE_OFN1040_n969), 
	.A(FE_OFN1039_n969));
   CLKBUFX2TS FE_OFC1039_n969 (.Y(FE_OFN1039_n969), 
	.A(n969));
   CLKBUFX2TS FE_OFC1038_n905 (.Y(FE_OFN1038_n905), 
	.A(FE_OFN1036_n905));
   CLKBUFX2TS FE_OFC1037_n905 (.Y(FE_OFN1037_n905), 
	.A(FE_OFN1034_n905));
   CLKBUFX2TS FE_OFC1036_n905 (.Y(FE_OFN1036_n905), 
	.A(FE_OFN1034_n905));
   CLKBUFX2TS FE_OFC1035_n905 (.Y(FE_OFN1035_n905), 
	.A(FE_OFN1034_n905));
   CLKBUFX2TS FE_OFC1034_n905 (.Y(FE_OFN1034_n905), 
	.A(n905));
   CLKBUFX2TS FE_OFC1033_n841 (.Y(FE_OFN1033_n841), 
	.A(FE_OFN1032_n841));
   CLKBUFX2TS FE_OFC1032_n841 (.Y(FE_OFN1032_n841), 
	.A(FE_OFN1031_n841));
   CLKBUFX2TS FE_OFC1031_n841 (.Y(FE_OFN1031_n841), 
	.A(FE_OFN1030_n841));
   CLKBUFX2TS FE_OFC1030_n841 (.Y(FE_OFN1030_n841), 
	.A(n841));
   CLKBUFX2TS FE_OFC1029_n777 (.Y(FE_OFN1029_n777), 
	.A(FE_OFN1027_n777));
   CLKBUFX2TS FE_OFC1028_n777 (.Y(FE_OFN1028_n777), 
	.A(FE_OFN1027_n777));
   CLKBUFX2TS FE_OFC1027_n777 (.Y(FE_OFN1027_n777), 
	.A(FE_OFN1026_n777));
   CLKBUFX2TS FE_OFC1026_n777 (.Y(FE_OFN1026_n777), 
	.A(n777));
   CLKBUFX2TS FE_OFC1025_n713 (.Y(FE_OFN1025_n713), 
	.A(FE_OFN1024_n713));
   CLKBUFX2TS FE_OFC1024_n713 (.Y(FE_OFN1024_n713), 
	.A(FE_OFN1023_n713));
   CLKBUFX2TS FE_OFC1023_n713 (.Y(FE_OFN1023_n713), 
	.A(FE_OFN1022_n713));
   CLKBUFX2TS FE_OFC1022_n713 (.Y(FE_OFN1022_n713), 
	.A(n713));
   CLKBUFX2TS FE_OFC1021_n649 (.Y(FE_OFN1021_n649), 
	.A(FE_OFN1020_n649));
   CLKBUFX2TS FE_OFC1020_n649 (.Y(FE_OFN1020_n649), 
	.A(FE_OFN1019_n649));
   CLKBUFX2TS FE_OFC1019_n649 (.Y(FE_OFN1019_n649), 
	.A(FE_OFN1018_n649));
   CLKBUFX2TS FE_OFC1018_n649 (.Y(FE_OFN1018_n649), 
	.A(n649));
   CLKBUFX2TS FE_OFC1017_n2569 (.Y(FE_OFN1017_n2569), 
	.A(FE_OFN1016_n2569));
   CLKBUFX2TS FE_OFC1016_n2569 (.Y(FE_OFN1016_n2569), 
	.A(FE_OFN1015_n2569));
   CLKBUFX2TS FE_OFC1015_n2569 (.Y(FE_OFN1015_n2569), 
	.A(FE_OFN1014_n2569));
   CLKBUFX2TS FE_OFC1014_n2569 (.Y(FE_OFN1014_n2569), 
	.A(n2569));
   CLKBUFX2TS FE_OFC1013_n1545 (.Y(FE_OFN1013_n1545), 
	.A(FE_OFN1012_n1545));
   CLKBUFX2TS FE_OFC1012_n1545 (.Y(FE_OFN1012_n1545), 
	.A(FE_OFN1010_n1545));
   CLKBUFX2TS FE_OFC1011_n1545 (.Y(FE_OFN1011_n1545), 
	.A(FE_OFN1010_n1545));
   CLKBUFX2TS FE_OFC1010_n1545 (.Y(FE_OFN1010_n1545), 
	.A(FE_OFN1009_n1545));
   CLKBUFX2TS FE_OFC1009_n1545 (.Y(FE_OFN1009_n1545), 
	.A(n1545));
   CLKBUFX2TS FE_OFC1008_n137 (.Y(FE_OFN1008_n137), 
	.A(FE_OFN1005_n137));
   CLKBUFX2TS FE_OFC1007_n137 (.Y(FE_OFN1007_n137), 
	.A(FE_OFN1006_n137));
   CLKBUFX2TS FE_OFC1006_n137 (.Y(FE_OFN1006_n137), 
	.A(FE_OFN1004_n137));
   CLKBUFX2TS FE_OFC1005_n137 (.Y(FE_OFN1005_n137), 
	.A(FE_OFN1004_n137));
   CLKBUFX2TS FE_OFC1004_n137 (.Y(FE_OFN1004_n137), 
	.A(n137));
   CLKBUFX2TS FE_OFC1003_n521 (.Y(FE_OFN1003_n521), 
	.A(FE_OFN1002_n521));
   CLKBUFX2TS FE_OFC1002_n521 (.Y(FE_OFN1002_n521), 
	.A(FE_OFN1001_n521));
   CLKBUFX2TS FE_OFC1001_n521 (.Y(FE_OFN1001_n521), 
	.A(FE_OFN1000_n521));
   CLKBUFX2TS FE_OFC1000_n521 (.Y(FE_OFN1000_n521), 
	.A(FE_OFN999_n521));
   CLKBUFX2TS FE_OFC999_n521 (.Y(FE_OFN999_n521), 
	.A(FE_OFN998_n521));
   CLKBUFX2TS FE_OFC998_n521 (.Y(FE_OFN998_n521), 
	.A(FE_OFN997_n521));
   CLKBUFX2TS FE_OFC997_n521 (.Y(FE_OFN997_n521), 
	.A(FE_OFN996_n521));
   CLKBUFX2TS FE_OFC996_n521 (.Y(FE_OFN996_n521), 
	.A(FE_OFN995_n521));
   CLKBUFX2TS FE_OFC995_n521 (.Y(FE_OFN995_n521), 
	.A(FE_OFN994_n521));
   CLKBUFX2TS FE_OFC994_n521 (.Y(FE_OFN994_n521), 
	.A(n521));
   CLKBUFX2TS FE_OFC993_n9431 (.Y(FE_OFN993_n9431), 
	.A(FE_OFN992_n9431));
   CLKBUFX2TS FE_OFC992_n9431 (.Y(FE_OFN992_n9431), 
	.A(FE_OFN991_n9431));
   CLKBUFX2TS FE_OFC991_n9431 (.Y(FE_OFN991_n9431), 
	.A(FE_OFN990_n9431));
   CLKBUFX2TS FE_OFC990_n9431 (.Y(FE_OFN990_n9431), 
	.A(FE_OFN988_n9431));
   CLKBUFX2TS FE_OFC989_n9431 (.Y(FE_OFN989_n9431), 
	.A(FE_OFN987_n9431));
   CLKBUFX2TS FE_OFC988_n9431 (.Y(FE_OFN988_n9431), 
	.A(FE_OFN986_n9431));
   CLKBUFX2TS FE_OFC987_n9431 (.Y(FE_OFN987_n9431), 
	.A(FE_OFN986_n9431));
   CLKBUFX2TS FE_OFC986_n9431 (.Y(FE_OFN986_n9431), 
	.A(FE_OFN985_n9431));
   CLKBUFX2TS FE_OFC985_n9431 (.Y(FE_OFN985_n9431), 
	.A(n9431));
   CLKBUFX2TS FE_OFC984_n9462 (.Y(FE_OFN984_n9462), 
	.A(FE_OFN983_n9462));
   CLKBUFX2TS FE_OFC983_n9462 (.Y(FE_OFN983_n9462), 
	.A(FE_OFN982_n9462));
   CLKBUFX2TS FE_OFC982_n9462 (.Y(FE_OFN982_n9462), 
	.A(FE_OFN981_n9462));
   CLKBUFX2TS FE_OFC981_n9462 (.Y(FE_OFN981_n9462), 
	.A(FE_OFN980_n9462));
   CLKBUFX2TS FE_OFC980_n9462 (.Y(FE_OFN980_n9462), 
	.A(FE_OFN978_n9462));
   CLKBUFX2TS FE_OFC979_n9462 (.Y(FE_OFN979_n9462), 
	.A(FE_OFN978_n9462));
   CLKBUFX2TS FE_OFC978_n9462 (.Y(FE_OFN978_n9462), 
	.A(FE_OFN977_n9462));
   CLKBUFX2TS FE_OFC977_n9462 (.Y(FE_OFN977_n9462), 
	.A(FE_OFN976_n9462));
   CLKBUFX2TS FE_OFC976_n9462 (.Y(FE_OFN976_n9462), 
	.A(FE_OFN974_n9462));
   CLKBUFX2TS FE_OFC975_n9462 (.Y(FE_OFN975_n9462), 
	.A(n9462));
   CLKBUFX2TS FE_OFC974_n9462 (.Y(FE_OFN974_n9462), 
	.A(n9462));
   CLKBUFX2TS FE_OFC973_n7207 (.Y(FE_OFN973_n7207), 
	.A(n7207));
   CLKBUFX2TS FE_OFC972_n3618 (.Y(FE_OFN972_n3618), 
	.A(FE_OFN971_n3618));
   CLKBUFX2TS FE_OFC971_n3618 (.Y(FE_OFN971_n3618), 
	.A(FE_OFN969_n3618));
   CLKBUFX2TS FE_OFC970_n3618 (.Y(FE_OFN970_n3618), 
	.A(FE_OFN969_n3618));
   CLKBUFX2TS FE_OFC969_n3618 (.Y(FE_OFN969_n3618), 
	.A(FE_OFN968_n3618));
   CLKBUFX2TS FE_OFC968_n3618 (.Y(FE_OFN968_n3618), 
	.A(FE_OFN967_n3618));
   CLKBUFX2TS FE_OFC967_n3618 (.Y(FE_OFN967_n3618), 
	.A(FE_OFN966_n3618));
   CLKBUFX2TS FE_OFC966_n3618 (.Y(FE_OFN966_n3618), 
	.A(FE_OFN965_n3618));
   CLKBUFX2TS FE_OFC965_n3618 (.Y(FE_OFN965_n3618), 
	.A(FE_OFN964_n3618));
   CLKBUFX2TS FE_OFC964_n3618 (.Y(FE_OFN964_n3618), 
	.A(FE_OFN962_n3618));
   CLKBUFX2TS FE_OFC963_n3618 (.Y(FE_OFN963_n3618), 
	.A(FE_OFN962_n3618));
   CLKBUFX2TS FE_OFC962_n3618 (.Y(FE_OFN962_n3618), 
	.A(n3618));
   CLKBUFX2TS FE_OFC961_n5467 (.Y(FE_OFN961_n5467), 
	.A(n5467));
   CLKBUFX2TS FE_OFC960_n3619 (.Y(FE_OFN960_n3619), 
	.A(FE_OFN959_n3619));
   CLKBUFX2TS FE_OFC959_n3619 (.Y(FE_OFN959_n3619), 
	.A(FE_OFN958_n3619));
   CLKBUFX2TS FE_OFC958_n3619 (.Y(FE_OFN958_n3619), 
	.A(FE_OFN957_n3619));
   CLKBUFX2TS FE_OFC957_n3619 (.Y(FE_OFN957_n3619), 
	.A(FE_OFN956_n3619));
   CLKBUFX2TS FE_OFC956_n3619 (.Y(FE_OFN956_n3619), 
	.A(FE_OFN955_n3619));
   CLKBUFX2TS FE_OFC955_n3619 (.Y(FE_OFN955_n3619), 
	.A(FE_OFN953_n3619));
   CLKBUFX2TS FE_OFC954_n3619 (.Y(FE_OFN954_n3619), 
	.A(FE_OFN952_n3619));
   CLKBUFX2TS FE_OFC953_n3619 (.Y(FE_OFN953_n3619), 
	.A(FE_OFN951_n3619));
   CLKBUFX2TS FE_OFC952_n3619 (.Y(FE_OFN952_n3619), 
	.A(FE_OFN951_n3619));
   CLKBUFX2TS FE_OFC951_n3619 (.Y(FE_OFN951_n3619), 
	.A(n3619));
   CLKBUFX2TS FE_OFC950_n3486 (.Y(FE_OFN950_n3486), 
	.A(FE_OFN949_n3486));
   CLKBUFX2TS FE_OFC949_n3486 (.Y(FE_OFN949_n3486), 
	.A(FE_OFN948_n3486));
   CLKBUFX2TS FE_OFC948_n3486 (.Y(FE_OFN948_n3486), 
	.A(FE_OFN947_n3486));
   CLKBUFX2TS FE_OFC947_n3486 (.Y(FE_OFN947_n3486), 
	.A(FE_OFN945_n3486));
   CLKBUFX2TS FE_OFC946_n3486 (.Y(FE_OFN946_n3486), 
	.A(FE_OFN944_n3486));
   CLKBUFX2TS FE_OFC945_n3486 (.Y(FE_OFN945_n3486), 
	.A(FE_OFN942_n3486));
   CLKBUFX2TS FE_OFC944_n3486 (.Y(FE_OFN944_n3486), 
	.A(FE_OFN943_n3486));
   CLKBUFX2TS FE_OFC943_n3486 (.Y(FE_OFN943_n3486), 
	.A(FE_OFN941_n3486));
   CLKBUFX2TS FE_OFC942_n3486 (.Y(FE_OFN942_n3486), 
	.A(FE_OFN940_n3486));
   CLKBUFX2TS FE_OFC941_n3486 (.Y(FE_OFN941_n3486), 
	.A(FE_OFN940_n3486));
   CLKBUFX2TS FE_OFC940_n3486 (.Y(FE_OFN940_n3486), 
	.A(n3486));
   CLKBUFX2TS FE_OFC939_n3487 (.Y(FE_OFN939_n3487), 
	.A(FE_OFN938_n3487));
   CLKBUFX2TS FE_OFC938_n3487 (.Y(FE_OFN938_n3487), 
	.A(FE_OFN937_n3487));
   CLKBUFX2TS FE_OFC937_n3487 (.Y(FE_OFN937_n3487), 
	.A(FE_OFN936_n3487));
   CLKBUFX2TS FE_OFC936_n3487 (.Y(FE_OFN936_n3487), 
	.A(FE_OFN935_n3487));
   CLKBUFX2TS FE_OFC935_n3487 (.Y(FE_OFN935_n3487), 
	.A(FE_OFN934_n3487));
   CLKBUFX2TS FE_OFC934_n3487 (.Y(FE_OFN934_n3487), 
	.A(FE_OFN932_n3487));
   CLKBUFX2TS FE_OFC933_n3487 (.Y(FE_OFN933_n3487), 
	.A(FE_OFN930_n3487));
   CLKBUFX2TS FE_OFC932_n3487 (.Y(FE_OFN932_n3487), 
	.A(FE_OFN931_n3487));
   CLKBUFX2TS FE_OFC931_n3487 (.Y(FE_OFN931_n3487), 
	.A(n3487));
   CLKBUFX2TS FE_OFC930_n3487 (.Y(FE_OFN930_n3487), 
	.A(n3487));
   CLKBUFX2TS FE_OFC929_n3574 (.Y(FE_OFN929_n3574), 
	.A(FE_OFN928_n3574));
   CLKBUFX2TS FE_OFC928_n3574 (.Y(FE_OFN928_n3574), 
	.A(FE_OFN927_n3574));
   CLKBUFX2TS FE_OFC927_n3574 (.Y(FE_OFN927_n3574), 
	.A(FE_OFN926_n3574));
   CLKBUFX2TS FE_OFC926_n3574 (.Y(FE_OFN926_n3574), 
	.A(FE_OFN925_n3574));
   CLKBUFX2TS FE_OFC925_n3574 (.Y(FE_OFN925_n3574), 
	.A(FE_OFN924_n3574));
   CLKBUFX2TS FE_OFC924_n3574 (.Y(FE_OFN924_n3574), 
	.A(FE_OFN923_n3574));
   CLKBUFX2TS FE_OFC923_n3574 (.Y(FE_OFN923_n3574), 
	.A(FE_OFN922_n3574));
   CLKBUFX2TS FE_OFC922_n3574 (.Y(FE_OFN922_n3574), 
	.A(FE_OFN920_n3574));
   CLKBUFX2TS FE_OFC921_n3574 (.Y(FE_OFN921_n3574), 
	.A(FE_OFN919_n3574));
   CLKBUFX2TS FE_OFC920_n3574 (.Y(FE_OFN920_n3574), 
	.A(FE_OFN919_n3574));
   CLKBUFX2TS FE_OFC919_n3574 (.Y(FE_OFN919_n3574), 
	.A(n3574));
   CLKBUFX2TS FE_OFC918_n3575 (.Y(FE_OFN918_n3575), 
	.A(FE_OFN917_n3575));
   CLKBUFX2TS FE_OFC917_n3575 (.Y(FE_OFN917_n3575), 
	.A(FE_OFN916_n3575));
   CLKBUFX2TS FE_OFC916_n3575 (.Y(FE_OFN916_n3575), 
	.A(FE_OFN915_n3575));
   CLKBUFX2TS FE_OFC915_n3575 (.Y(FE_OFN915_n3575), 
	.A(FE_OFN914_n3575));
   CLKBUFX2TS FE_OFC914_n3575 (.Y(FE_OFN914_n3575), 
	.A(FE_OFN913_n3575));
   CLKBUFX2TS FE_OFC913_n3575 (.Y(FE_OFN913_n3575), 
	.A(FE_OFN912_n3575));
   CLKBUFX2TS FE_OFC912_n3575 (.Y(FE_OFN912_n3575), 
	.A(FE_OFN911_n3575));
   CLKBUFX2TS FE_OFC911_n3575 (.Y(FE_OFN911_n3575), 
	.A(FE_OFN910_n3575));
   CLKBUFX2TS FE_OFC910_n3575 (.Y(FE_OFN910_n3575), 
	.A(FE_OFN909_n3575));
   CLKBUFX2TS FE_OFC909_n3575 (.Y(FE_OFN909_n3575), 
	.A(n3575));
   CLKBUFX2TS FE_OFC908_n3530 (.Y(FE_OFN908_n3530), 
	.A(FE_OFN905_n3530));
   CLKBUFX2TS FE_OFC907_n3530 (.Y(FE_OFN907_n3530), 
	.A(FE_OFN904_n3530));
   CLKBUFX2TS FE_OFC906_n3530 (.Y(FE_OFN906_n3530), 
	.A(FE_OFN904_n3530));
   CLKBUFX2TS FE_OFC905_n3530 (.Y(FE_OFN905_n3530), 
	.A(FE_OFN902_n3530));
   CLKBUFX2TS FE_OFC904_n3530 (.Y(FE_OFN904_n3530), 
	.A(FE_OFN903_n3530));
   CLKBUFX2TS FE_OFC903_n3530 (.Y(FE_OFN903_n3530), 
	.A(FE_OFN901_n3530));
   CLKBUFX2TS FE_OFC902_n3530 (.Y(FE_OFN902_n3530), 
	.A(FE_OFN901_n3530));
   CLKBUFX2TS FE_OFC901_n3530 (.Y(FE_OFN901_n3530), 
	.A(FE_OFN899_n3530));
   CLKBUFX2TS FE_OFC900_n3530 (.Y(FE_OFN900_n3530), 
	.A(FE_OFN899_n3530));
   CLKBUFX2TS FE_OFC899_n3530 (.Y(FE_OFN899_n3530), 
	.A(FE_OFN898_n3530));
   CLKBUFX2TS FE_OFC898_n3530 (.Y(FE_OFN898_n3530), 
	.A(n3530));
   CLKBUFX2TS FE_OFC897_n3531 (.Y(FE_OFN897_n3531), 
	.A(FE_OFN894_n3531));
   CLKBUFX2TS FE_OFC896_n3531 (.Y(FE_OFN896_n3531), 
	.A(FE_OFN895_n3531));
   CLKBUFX2TS FE_OFC895_n3531 (.Y(FE_OFN895_n3531), 
	.A(FE_OFN891_n3531));
   CLKBUFX2TS FE_OFC894_n3531 (.Y(FE_OFN894_n3531), 
	.A(FE_OFN893_n3531));
   CLKBUFX2TS FE_OFC893_n3531 (.Y(FE_OFN893_n3531), 
	.A(FE_OFN888_n3531));
   CLKBUFX2TS FE_OFC892_n3531 (.Y(FE_OFN892_n3531), 
	.A(FE_OFN889_n3531));
   CLKBUFX2TS FE_OFC891_n3531 (.Y(FE_OFN891_n3531), 
	.A(FE_OFN888_n3531));
   CLKBUFX2TS FE_OFC890_n3531 (.Y(FE_OFN890_n3531), 
	.A(FE_OFN889_n3531));
   CLKBUFX2TS FE_OFC889_n3531 (.Y(FE_OFN889_n3531), 
	.A(n3531));
   CLKBUFX2TS FE_OFC888_n3531 (.Y(FE_OFN888_n3531), 
	.A(n3531));
   CLKBUFX2TS FE_OFC887_n3662 (.Y(FE_OFN887_n3662), 
	.A(FE_OFN885_n3662));
   CLKBUFX2TS FE_OFC886_n3662 (.Y(FE_OFN886_n3662), 
	.A(FE_OFN884_n3662));
   CLKBUFX2TS FE_OFC885_n3662 (.Y(FE_OFN885_n3662), 
	.A(FE_OFN882_n3662));
   CLKBUFX2TS FE_OFC884_n3662 (.Y(FE_OFN884_n3662), 
	.A(FE_OFN883_n3662));
   CLKBUFX2TS FE_OFC883_n3662 (.Y(FE_OFN883_n3662), 
	.A(FE_OFN880_n3662));
   CLKBUFX2TS FE_OFC882_n3662 (.Y(FE_OFN882_n3662), 
	.A(FE_OFN881_n3662));
   CLKBUFX2TS FE_OFC881_n3662 (.Y(FE_OFN881_n3662), 
	.A(FE_OFN880_n3662));
   CLKBUFX2TS FE_OFC880_n3662 (.Y(FE_OFN880_n3662), 
	.A(FE_OFN879_n3662));
   CLKBUFX2TS FE_OFC879_n3662 (.Y(FE_OFN879_n3662), 
	.A(FE_OFN878_n3662));
   CLKBUFX2TS FE_OFC878_n3662 (.Y(FE_OFN878_n3662), 
	.A(FE_OFN877_n3662));
   CLKBUFX2TS FE_OFC877_n3662 (.Y(FE_OFN877_n3662), 
	.A(n3662));
   CLKBUFX2TS FE_OFC876_n3663 (.Y(FE_OFN876_n3663), 
	.A(FE_OFN874_n3663));
   CLKBUFX2TS FE_OFC875_n3663 (.Y(FE_OFN875_n3663), 
	.A(FE_OFN873_n3663));
   CLKBUFX2TS FE_OFC874_n3663 (.Y(FE_OFN874_n3663), 
	.A(FE_OFN872_n3663));
   CLKBUFX2TS FE_OFC873_n3663 (.Y(FE_OFN873_n3663), 
	.A(FE_OFN870_n3663));
   CLKBUFX2TS FE_OFC872_n3663 (.Y(FE_OFN872_n3663), 
	.A(FE_OFN870_n3663));
   CLKBUFX2TS FE_OFC871_n3663 (.Y(FE_OFN871_n3663), 
	.A(FE_OFN869_n3663));
   CLKBUFX2TS FE_OFC870_n3663 (.Y(FE_OFN870_n3663), 
	.A(FE_OFN868_n3663));
   CLKBUFX2TS FE_OFC869_n3663 (.Y(FE_OFN869_n3663), 
	.A(FE_OFN867_n3663));
   CLKBUFX2TS FE_OFC868_n3663 (.Y(FE_OFN868_n3663), 
	.A(n3663));
   CLKBUFX2TS FE_OFC867_n3663 (.Y(FE_OFN867_n3663), 
	.A(n3663));
   CLKBUFX2TS FE_OFC866_n7015 (.Y(FE_OFN866_n7015), 
	.A(FE_OFN865_n7015));
   CLKBUFX2TS FE_OFC865_n7015 (.Y(FE_OFN865_n7015), 
	.A(FE_OFN863_n7015));
   CLKBUFX2TS FE_OFC864_n7015 (.Y(FE_OFN864_n7015), 
	.A(FE_OFN862_n7015));
   CLKBUFX2TS FE_OFC863_n7015 (.Y(FE_OFN863_n7015), 
	.A(FE_OFN862_n7015));
   CLKBUFX2TS FE_OFC862_n7015 (.Y(FE_OFN862_n7015), 
	.A(n7015));
   CLKBUFX2TS FE_OFC861_n7017 (.Y(FE_OFN861_n7017), 
	.A(FE_OFN860_n7017));
   CLKBUFX2TS FE_OFC860_n7017 (.Y(FE_OFN860_n7017), 
	.A(FE_OFN859_n7017));
   CLKBUFX2TS FE_OFC859_n7017 (.Y(FE_OFN859_n7017), 
	.A(FE_OFN858_n7017));
   CLKBUFX2TS FE_OFC858_n7017 (.Y(FE_OFN858_n7017), 
	.A(FE_OFN857_n7017));
   CLKBUFX2TS FE_OFC857_n7017 (.Y(FE_OFN857_n7017), 
	.A(n7017));
   CLKBUFX2TS FE_OFC856_n7018 (.Y(FE_OFN856_n7018), 
	.A(FE_OFN855_n7018));
   CLKBUFX2TS FE_OFC855_n7018 (.Y(FE_OFN855_n7018), 
	.A(FE_OFN853_n7018));
   CLKBUFX2TS FE_OFC854_n7018 (.Y(FE_OFN854_n7018), 
	.A(FE_OFN853_n7018));
   CLKBUFX2TS FE_OFC853_n7018 (.Y(FE_OFN853_n7018), 
	.A(n7018));
   CLKBUFX2TS FE_OFC852_n7016 (.Y(FE_OFN852_n7016), 
	.A(FE_OFN851_n7016));
   CLKBUFX2TS FE_OFC851_n7016 (.Y(FE_OFN851_n7016), 
	.A(FE_OFN850_n7016));
   CLKBUFX2TS FE_OFC850_n7016 (.Y(FE_OFN850_n7016), 
	.A(FE_OFN849_n7016));
   CLKBUFX2TS FE_OFC849_n7016 (.Y(FE_OFN849_n7016), 
	.A(n7016));
   CLKBUFX3TS FE_OFC848_ram_write_enable (.Y(ram_write_enable), 
	.A(FE_OFN848_ram_write_enable));
   CLKBUFX2TS FE_OFC847_n7619 (.Y(FE_OFN847_n7619), 
	.A(FE_OFN844_n7619));
   CLKBUFX2TS FE_OFC846_n7619 (.Y(FE_OFN846_n7619), 
	.A(FE_OFN845_n7619));
   CLKBUFX2TS FE_OFC845_n7619 (.Y(FE_OFN845_n7619), 
	.A(FE_OFN841_n7619));
   CLKBUFX2TS FE_OFC844_n7619 (.Y(FE_OFN844_n7619), 
	.A(FE_OFN840_n7619));
   CLKBUFX2TS FE_OFC843_n7619 (.Y(FE_OFN843_n7619), 
	.A(FE_OFN839_n7619));
   CLKBUFX2TS FE_OFC842_n7619 (.Y(FE_OFN842_n7619), 
	.A(FE_OFN838_n7619));
   CLKBUFX2TS FE_OFC841_n7619 (.Y(FE_OFN841_n7619), 
	.A(FE_OFN837_n7619));
   CLKBUFX2TS FE_OFC840_n7619 (.Y(FE_OFN840_n7619), 
	.A(FE_OFN836_n7619));
   CLKBUFX2TS FE_OFC839_n7619 (.Y(FE_OFN839_n7619), 
	.A(FE_OFN833_n7619));
   CLKBUFX2TS FE_OFC838_n7619 (.Y(FE_OFN838_n7619), 
	.A(FE_OFN834_n7619));
   CLKBUFX2TS FE_OFC837_n7619 (.Y(FE_OFN837_n7619), 
	.A(FE_OFN831_n7619));
   CLKBUFX2TS FE_OFC836_n7619 (.Y(FE_OFN836_n7619), 
	.A(FE_OFN830_n7619));
   CLKBUFX2TS FE_OFC835_n7619 (.Y(FE_OFN835_n7619), 
	.A(FE_OFN832_n7619));
   CLKBUFX2TS FE_OFC834_n7619 (.Y(FE_OFN834_n7619), 
	.A(FE_OFN826_n7619));
   CLKBUFX2TS FE_OFC833_n7619 (.Y(FE_OFN833_n7619), 
	.A(FE_OFN828_n7619));
   CLKBUFX2TS FE_OFC832_n7619 (.Y(FE_OFN832_n7619), 
	.A(FE_OFN825_n7619));
   CLKBUFX2TS FE_OFC831_n7619 (.Y(FE_OFN831_n7619), 
	.A(FE_OFN822_n7619));
   CLKBUFX2TS FE_OFC830_n7619 (.Y(FE_OFN830_n7619), 
	.A(FE_OFN824_n7619));
   CLKBUFX2TS FE_OFC829_n7619 (.Y(FE_OFN829_n7619), 
	.A(FE_OFN822_n7619));
   CLKBUFX2TS FE_OFC828_n7619 (.Y(FE_OFN828_n7619), 
	.A(FE_OFN821_n7619));
   CLKBUFX2TS FE_OFC827_n7619 (.Y(FE_OFN827_n7619), 
	.A(FE_OFN824_n7619));
   CLKBUFX2TS FE_OFC826_n7619 (.Y(FE_OFN826_n7619), 
	.A(FE_OFN819_n7619));
   CLKBUFX2TS FE_OFC825_n7619 (.Y(FE_OFN825_n7619), 
	.A(FE_OFN818_n7619));
   CLKBUFX2TS FE_OFC824_n7619 (.Y(FE_OFN824_n7619), 
	.A(FE_OFN820_n7619));
   CLKBUFX2TS FE_OFC823_n7619 (.Y(FE_OFN823_n7619), 
	.A(FE_OFN816_n7619));
   CLKBUFX2TS FE_OFC822_n7619 (.Y(FE_OFN822_n7619), 
	.A(FE_OFN817_n7619));
   CLKBUFX2TS FE_OFC821_n7619 (.Y(FE_OFN821_n7619), 
	.A(FE_OFN809_n7619));
   CLKBUFX2TS FE_OFC820_n7619 (.Y(FE_OFN820_n7619), 
	.A(FE_OFN813_n7619));
   CLKBUFX2TS FE_OFC819_n7619 (.Y(FE_OFN819_n7619), 
	.A(FE_OFN814_n7619));
   CLKBUFX2TS FE_OFC818_n7619 (.Y(FE_OFN818_n7619), 
	.A(FE_OFN812_n7619));
   CLKBUFX2TS FE_OFC817_n7619 (.Y(FE_OFN817_n7619), 
	.A(FE_OFN812_n7619));
   CLKBUFX2TS FE_OFC816_n7619 (.Y(FE_OFN816_n7619), 
	.A(FE_OFN810_n7619));
   CLKBUFX2TS FE_OFC815_n7619 (.Y(FE_OFN815_n7619), 
	.A(FE_OFN808_n7619));
   CLKBUFX2TS FE_OFC814_n7619 (.Y(FE_OFN814_n7619), 
	.A(FE_OFN810_n7619));
   CLKBUFX2TS FE_OFC813_n7619 (.Y(FE_OFN813_n7619), 
	.A(FE_OFN806_n7619));
   CLKBUFX2TS FE_OFC812_n7619 (.Y(FE_OFN812_n7619), 
	.A(FE_OFN803_n7619));
   CLKBUFX2TS FE_OFC811_n7619 (.Y(FE_OFN811_n7619), 
	.A(FE_OFN804_n7619));
   CLKBUFX2TS FE_OFC810_n7619 (.Y(FE_OFN810_n7619), 
	.A(FE_OFN805_n7619));
   CLKBUFX2TS FE_OFC809_n7619 (.Y(FE_OFN809_n7619), 
	.A(FE_OFN804_n7619));
   CLKBUFX2TS FE_OFC808_n7619 (.Y(FE_OFN808_n7619), 
	.A(FE_OFN803_n7619));
   CLKBUFX2TS FE_OFC807_n7619 (.Y(FE_OFN807_n7619), 
	.A(FE_OFN803_n7619));
   CLKBUFX2TS FE_OFC806_n7619 (.Y(FE_OFN806_n7619), 
	.A(FE_OFN801_n7619));
   CLKBUFX2TS FE_OFC805_n7619 (.Y(FE_OFN805_n7619), 
	.A(FE_OFN798_n7619));
   CLKBUFX2TS FE_OFC804_n7619 (.Y(FE_OFN804_n7619), 
	.A(FE_OFN799_n7619));
   CLKBUFX2TS FE_OFC803_n7619 (.Y(FE_OFN803_n7619), 
	.A(FE_OFN795_n7619));
   CLKBUFX2TS FE_OFC802_n7619 (.Y(FE_OFN802_n7619), 
	.A(FE_OFN796_n7619));
   CLKBUFX2TS FE_OFC801_n7619 (.Y(FE_OFN801_n7619), 
	.A(FE_OFN796_n7619));
   CLKBUFX2TS FE_OFC800_n7619 (.Y(FE_OFN800_n7619), 
	.A(FE_OFN790_n7619));
   CLKBUFX2TS FE_OFC799_n7619 (.Y(FE_OFN799_n7619), 
	.A(FE_OFN793_n7619));
   CLKBUFX2TS FE_OFC798_n7619 (.Y(FE_OFN798_n7619), 
	.A(FE_OFN794_n7619));
   CLKBUFX2TS FE_OFC797_n7619 (.Y(FE_OFN797_n7619), 
	.A(FE_OFN794_n7619));
   CLKBUFX2TS FE_OFC796_n7619 (.Y(FE_OFN796_n7619), 
	.A(FE_OFN792_n7619));
   CLKBUFX2TS FE_OFC795_n7619 (.Y(FE_OFN795_n7619), 
	.A(FE_OFN791_n7619));
   CLKBUFX2TS FE_OFC794_n7619 (.Y(FE_OFN794_n7619), 
	.A(FE_OFN792_n7619));
   CLKBUFX2TS FE_OFC793_n7619 (.Y(FE_OFN793_n7619), 
	.A(FE_OFN788_n7619));
   CLKBUFX2TS FE_OFC792_n7619 (.Y(FE_OFN792_n7619), 
	.A(FE_OFN786_n7619));
   CLKBUFX2TS FE_OFC791_n7619 (.Y(FE_OFN791_n7619), 
	.A(FE_OFN789_n7619));
   CLKBUFX2TS FE_OFC790_n7619 (.Y(FE_OFN790_n7619), 
	.A(FE_OFN787_n7619));
   CLKBUFX2TS FE_OFC789_n7619 (.Y(FE_OFN789_n7619), 
	.A(FE_OFN785_n7619));
   CLKBUFX2TS FE_OFC788_n7619 (.Y(FE_OFN788_n7619), 
	.A(FE_OFN784_n7619));
   CLKBUFX2TS FE_OFC787_n7619 (.Y(FE_OFN787_n7619), 
	.A(FE_OFN782_n7619));
   CLKBUFX2TS FE_OFC786_n7619 (.Y(FE_OFN786_n7619), 
	.A(FE_OFN783_n7619));
   CLKBUFX2TS FE_OFC785_n7619 (.Y(FE_OFN785_n7619), 
	.A(FE_OFN781_n7619));
   CLKBUFX2TS FE_OFC784_n7619 (.Y(FE_OFN784_n7619), 
	.A(FE_OFN781_n7619));
   CLKBUFX2TS FE_OFC783_n7619 (.Y(FE_OFN783_n7619), 
	.A(FE_OFN780_n7619));
   CLKBUFX2TS FE_OFC782_n7619 (.Y(FE_OFN782_n7619), 
	.A(FE_OFN780_n7619));
   CLKBUFX2TS FE_OFC781_n7619 (.Y(FE_OFN781_n7619), 
	.A(FE_OFN777_n7619));
   CLKBUFX2TS FE_OFC780_n7619 (.Y(FE_OFN780_n7619), 
	.A(FE_OFN778_n7619));
   CLKBUFX2TS FE_OFC779_n7619 (.Y(FE_OFN779_n7619), 
	.A(FE_OFN778_n7619));
   CLKBUFX2TS FE_OFC778_n7619 (.Y(FE_OFN778_n7619), 
	.A(n7619));
   CLKBUFX2TS FE_OFC777_n7619 (.Y(FE_OFN777_n7619), 
	.A(n7619));
   CLKBUFX2TS FE_OFC776_n3829 (.Y(FE_OFN776_n3829), 
	.A(n3829));
   CLKBUFX2TS FE_OFC775_n3720 (.Y(FE_OFN775_n3720), 
	.A(FE_OFN774_n3720));
   CLKBUFX2TS FE_OFC774_n3720 (.Y(FE_OFN774_n3720), 
	.A(FE_OFN772_n3720));
   CLKBUFX2TS FE_OFC773_n3720 (.Y(FE_OFN773_n3720), 
	.A(FE_OFN772_n3720));
   CLKBUFX2TS FE_OFC772_n3720 (.Y(FE_OFN772_n3720), 
	.A(FE_OFN771_n3720));
   CLKBUFX2TS FE_OFC771_n3720 (.Y(FE_OFN771_n3720), 
	.A(FE_OFN769_n3720));
   CLKBUFX2TS FE_OFC770_n3720 (.Y(FE_OFN770_n3720), 
	.A(FE_OFN769_n3720));
   CLKBUFX2TS FE_OFC769_n3720 (.Y(FE_OFN769_n3720), 
	.A(FE_OFN768_n3720));
   CLKBUFX2TS FE_OFC768_n3720 (.Y(FE_OFN768_n3720), 
	.A(FE_OFN766_n3720));
   CLKBUFX2TS FE_OFC767_n3720 (.Y(FE_OFN767_n3720), 
	.A(FE_OFN765_n3720));
   CLKBUFX2TS FE_OFC766_n3720 (.Y(FE_OFN766_n3720), 
	.A(FE_OFN765_n3720));
   CLKBUFX2TS FE_OFC765_n3720 (.Y(FE_OFN765_n3720), 
	.A(n3720));
   CLKBUFX2TS FE_OFC764_n3721 (.Y(FE_OFN764_n3721), 
	.A(FE_OFN763_n3721));
   CLKBUFX2TS FE_OFC763_n3721 (.Y(FE_OFN763_n3721), 
	.A(FE_OFN761_n3721));
   CLKBUFX2TS FE_OFC762_n3721 (.Y(FE_OFN762_n3721), 
	.A(FE_OFN761_n3721));
   CLKBUFX2TS FE_OFC761_n3721 (.Y(FE_OFN761_n3721), 
	.A(FE_OFN760_n3721));
   CLKBUFX2TS FE_OFC760_n3721 (.Y(FE_OFN760_n3721), 
	.A(FE_OFN758_n3721));
   CLKBUFX2TS FE_OFC759_n3721 (.Y(FE_OFN759_n3721), 
	.A(FE_OFN758_n3721));
   CLKBUFX2TS FE_OFC758_n3721 (.Y(FE_OFN758_n3721), 
	.A(FE_OFN757_n3721));
   CLKBUFX2TS FE_OFC757_n3721 (.Y(FE_OFN757_n3721), 
	.A(FE_OFN756_n3721));
   CLKBUFX2TS FE_OFC756_n3721 (.Y(FE_OFN756_n3721), 
	.A(n3721));
   CLKBUFX2TS FE_OFC755_n3721 (.Y(FE_OFN755_n3721), 
	.A(n3721));
   CLKBUFX2TS FE_OFC754_n3722 (.Y(FE_OFN754_n3722), 
	.A(FE_OFN753_n3722));
   CLKBUFX2TS FE_OFC753_n3722 (.Y(FE_OFN753_n3722), 
	.A(FE_OFN751_n3722));
   CLKBUFX2TS FE_OFC752_n3722 (.Y(FE_OFN752_n3722), 
	.A(FE_OFN751_n3722));
   CLKBUFX2TS FE_OFC751_n3722 (.Y(FE_OFN751_n3722), 
	.A(FE_OFN750_n3722));
   CLKBUFX2TS FE_OFC750_n3722 (.Y(FE_OFN750_n3722), 
	.A(FE_OFN748_n3722));
   CLKBUFX2TS FE_OFC749_n3722 (.Y(FE_OFN749_n3722), 
	.A(FE_OFN748_n3722));
   CLKBUFX2TS FE_OFC748_n3722 (.Y(FE_OFN748_n3722), 
	.A(FE_OFN747_n3722));
   CLKBUFX2TS FE_OFC747_n3722 (.Y(FE_OFN747_n3722), 
	.A(FE_OFN745_n3722));
   CLKBUFX2TS FE_OFC746_n3722 (.Y(FE_OFN746_n3722), 
	.A(n3722));
   CLKBUFX2TS FE_OFC745_n3722 (.Y(FE_OFN745_n3722), 
	.A(n3722));
   CLKBUFX2TS FE_OFC744_n4829 (.Y(FE_OFN744_n4829), 
	.A(FE_OFN743_n4829));
   CLKBUFX2TS FE_OFC743_n4829 (.Y(FE_OFN743_n4829), 
	.A(FE_OFN740_n4829));
   CLKBUFX2TS FE_OFC742_n4829 (.Y(FE_OFN742_n4829), 
	.A(FE_OFN741_n4829));
   CLKBUFX2TS FE_OFC741_n4829 (.Y(FE_OFN741_n4829), 
	.A(FE_OFN739_n4829));
   CLKBUFX2TS FE_OFC740_n4829 (.Y(FE_OFN740_n4829), 
	.A(FE_OFN738_n4829));
   CLKBUFX2TS FE_OFC739_n4829 (.Y(FE_OFN739_n4829), 
	.A(FE_OFN737_n4829));
   CLKBUFX2TS FE_OFC738_n4829 (.Y(FE_OFN738_n4829), 
	.A(FE_OFN737_n4829));
   CLKBUFX2TS FE_OFC737_n4829 (.Y(FE_OFN737_n4829), 
	.A(FE_OFN736_n4829));
   CLKBUFX2TS FE_OFC736_n4829 (.Y(FE_OFN736_n4829), 
	.A(n4829));
   CLKBUFX2TS FE_OFC735_n4829 (.Y(FE_OFN735_n4829), 
	.A(n4829));
   CLKBUFX2TS FE_OFC734_n8057 (.Y(FE_OFN734_n8057), 
	.A(FE_OFN733_n8057));
   CLKBUFX2TS FE_OFC733_n8057 (.Y(FE_OFN733_n8057), 
	.A(FE_OFN732_n8057));
   CLKBUFX2TS FE_OFC732_n8057 (.Y(FE_OFN732_n8057), 
	.A(n8057));
   CLKBUFX2TS FE_OFC731_n8058 (.Y(FE_OFN731_n8058), 
	.A(FE_OFN730_n8058));
   CLKBUFX2TS FE_OFC730_n8058 (.Y(FE_OFN730_n8058), 
	.A(FE_OFN729_n8058));
   CLKBUFX2TS FE_OFC729_n8058 (.Y(FE_OFN729_n8058), 
	.A(n8058));
   CLKBUFX2TS FE_OFC728_n4643 (.Y(FE_OFN728_n4643), 
	.A(FE_OFN727_n4643));
   CLKBUFX2TS FE_OFC727_n4643 (.Y(FE_OFN727_n4643), 
	.A(FE_OFN725_n4643));
   CLKBUFX2TS FE_OFC726_n4643 (.Y(FE_OFN726_n4643), 
	.A(FE_OFN725_n4643));
   CLKBUFX2TS FE_OFC725_n4643 (.Y(FE_OFN725_n4643), 
	.A(FE_OFN724_n4643));
   CLKBUFX2TS FE_OFC724_n4643 (.Y(FE_OFN724_n4643), 
	.A(FE_OFN723_n4643));
   CLKBUFX2TS FE_OFC723_n4643 (.Y(FE_OFN723_n4643), 
	.A(FE_OFN722_n4643));
   CLKBUFX2TS FE_OFC722_n4643 (.Y(FE_OFN722_n4643), 
	.A(FE_OFN720_n4643));
   CLKBUFX2TS FE_OFC721_n4643 (.Y(FE_OFN721_n4643), 
	.A(FE_OFN1823_n4643));
   CLKBUFX2TS FE_OFC720_n4643 (.Y(FE_OFN720_n4643), 
	.A(FE_OFN1823_n4643));
   CLKBUFX2TS FE_OFC719_n4643 (.Y(FE_OFN719_n4643), 
	.A(n4643));
   CLKBUFX2TS FE_OFC718_n8051 (.Y(FE_OFN718_n8051), 
	.A(FE_OFN717_n8051));
   CLKBUFX2TS FE_OFC717_n8051 (.Y(FE_OFN717_n8051), 
	.A(n8051));
   CLKBUFX2TS FE_OFC716_n4207 (.Y(FE_OFN716_n4207), 
	.A(FE_OFN714_n4207));
   CLKBUFX2TS FE_OFC715_n4207 (.Y(FE_OFN715_n4207), 
	.A(FE_OFN712_n4207));
   CLKBUFX2TS FE_OFC714_n4207 (.Y(FE_OFN714_n4207), 
	.A(FE_OFN712_n4207));
   CLKBUFX2TS FE_OFC713_n4207 (.Y(FE_OFN713_n4207), 
	.A(FE_OFN710_n4207));
   CLKBUFX2TS FE_OFC712_n4207 (.Y(FE_OFN712_n4207), 
	.A(FE_OFN710_n4207));
   CLKBUFX2TS FE_OFC711_n4207 (.Y(FE_OFN711_n4207), 
	.A(FE_OFN709_n4207));
   CLKBUFX2TS FE_OFC710_n4207 (.Y(FE_OFN710_n4207), 
	.A(FE_OFN709_n4207));
   CLKBUFX2TS FE_OFC709_n4207 (.Y(FE_OFN709_n4207), 
	.A(n4207));
   CLKBUFX2TS FE_OFC708_n3959 (.Y(FE_OFN708_n3959), 
	.A(FE_OFN705_n3959));
   CLKBUFX2TS FE_OFC707_n3959 (.Y(FE_OFN707_n3959), 
	.A(FE_OFN703_n3959));
   CLKBUFX2TS FE_OFC706_n3959 (.Y(FE_OFN706_n3959), 
	.A(FE_OFN703_n3959));
   CLKBUFX2TS FE_OFC705_n3959 (.Y(FE_OFN705_n3959), 
	.A(FE_OFN702_n3959));
   CLKBUFX2TS FE_OFC704_n3959 (.Y(FE_OFN704_n3959), 
	.A(FE_OFN701_n3959));
   CLKBUFX2TS FE_OFC703_n3959 (.Y(FE_OFN703_n3959), 
	.A(FE_OFN702_n3959));
   CLKBUFX2TS FE_OFC702_n3959 (.Y(FE_OFN702_n3959), 
	.A(FE_OFN699_n3959));
   CLKBUFX2TS FE_OFC701_n3959 (.Y(FE_OFN701_n3959), 
	.A(FE_OFN699_n3959));
   CLKBUFX2TS FE_OFC700_n3959 (.Y(FE_OFN700_n3959), 
	.A(n3959));
   CLKBUFX2TS FE_OFC699_n3959 (.Y(FE_OFN699_n3959), 
	.A(n3959));
   CLKBUFX2TS FE_OFC698_n8052 (.Y(FE_OFN698_n8052), 
	.A(FE_OFN696_n8052));
   CLKBUFX2TS FE_OFC697_n8052 (.Y(FE_OFN697_n8052), 
	.A(FE_OFN696_n8052));
   CLKBUFX2TS FE_OFC696_n8052 (.Y(FE_OFN696_n8052), 
	.A(n8052));
   CLKBUFX2TS FE_OFC695_n4134 (.Y(FE_OFN695_n4134), 
	.A(FE_OFN694_n4134));
   CLKBUFX2TS FE_OFC694_n4134 (.Y(FE_OFN694_n4134), 
	.A(FE_OFN693_n4134));
   CLKINVX1TS FE_OFC693_n4134 (.Y(FE_OFN693_n4134), 
	.A(FE_OFN690_n4134));
   CLKINVX1TS FE_OFC692_n4134 (.Y(FE_OFN692_n4134), 
	.A(FE_OFN690_n4134));
   CLKINVX1TS FE_OFC691_n4134 (.Y(FE_OFN691_n4134), 
	.A(FE_OFN690_n4134));
   CLKINVX1TS FE_OFC690_n4134 (.Y(FE_OFN690_n4134), 
	.A(FE_OFN689_n4134));
   CLKBUFX2TS FE_OFC689_n4134 (.Y(FE_OFN689_n4134), 
	.A(FE_OFN688_n4134));
   CLKBUFX2TS FE_OFC688_n4134 (.Y(FE_OFN688_n4134), 
	.A(FE_OFN687_n4134));
   CLKBUFX2TS FE_OFC687_n4134 (.Y(FE_OFN687_n4134), 
	.A(FE_OFN685_n4134));
   CLKBUFX2TS FE_OFC686_n4134 (.Y(FE_OFN686_n4134), 
	.A(FE_OFN685_n4134));
   CLKBUFX2TS FE_OFC685_n4134 (.Y(FE_OFN685_n4134), 
	.A(FE_OFN684_n4134));
   CLKBUFX2TS FE_OFC684_n4134 (.Y(FE_OFN684_n4134), 
	.A(FE_OFN683_n4134));
   CLKBUFX2TS FE_OFC683_n4134 (.Y(FE_OFN683_n4134), 
	.A(n4134));
   CLKBUFX2TS FE_OFC682_n8050 (.Y(FE_OFN682_n8050), 
	.A(FE_OFN681_n8050));
   CLKBUFX2TS FE_OFC681_n8050 (.Y(FE_OFN681_n8050), 
	.A(FE_OFN680_n8050));
   CLKBUFX2TS FE_OFC680_n8050 (.Y(FE_OFN680_n8050), 
	.A(n8050));
   CLKBUFX2TS FE_OFC679_n8050 (.Y(FE_OFN679_n8050), 
	.A(n8050));
   CLKBUFX2TS FE_OFC678_n7295 (.Y(FE_OFN678_n7295), 
	.A(n7295));
   CLKBUFX2TS FE_OFC677_n4759 (.Y(FE_OFN677_n4759), 
	.A(FE_OFN676_n4759));
   CLKBUFX2TS FE_OFC676_n4759 (.Y(FE_OFN676_n4759), 
	.A(FE_OFN674_n4759));
   CLKBUFX2TS FE_OFC675_n4759 (.Y(FE_OFN675_n4759), 
	.A(FE_OFN674_n4759));
   CLKBUFX2TS FE_OFC674_n4759 (.Y(FE_OFN674_n4759), 
	.A(FE_OFN673_n4759));
   CLKBUFX2TS FE_OFC673_n4759 (.Y(FE_OFN673_n4759), 
	.A(FE_OFN672_n4759));
   CLKBUFX2TS FE_OFC672_n4759 (.Y(FE_OFN672_n4759), 
	.A(FE_OFN671_n4759));
   CLKBUFX2TS FE_OFC671_n4759 (.Y(FE_OFN671_n4759), 
	.A(FE_OFN670_n4759));
   CLKBUFX2TS FE_OFC670_n4759 (.Y(FE_OFN670_n4759), 
	.A(FE_OFN668_n4759));
   CLKBUFX2TS FE_OFC669_n4759 (.Y(FE_OFN669_n4759), 
	.A(FE_OFN667_n4759));
   CLKBUFX2TS FE_OFC668_n4759 (.Y(FE_OFN668_n4759), 
	.A(FE_OFN667_n4759));
   CLKBUFX2TS FE_OFC667_n4759 (.Y(FE_OFN667_n4759), 
	.A(FE_OFN666_n4759));
   CLKBUFX2TS FE_OFC666_n4759 (.Y(FE_OFN666_n4759), 
	.A(n4759));
   CLKBUFX2TS FE_OFC665_n8053 (.Y(FE_OFN665_n8053), 
	.A(FE_OFN664_n8053));
   CLKBUFX2TS FE_OFC664_n8053 (.Y(FE_OFN664_n8053), 
	.A(n8053));
   CLKBUFX2TS FE_OFC663_n4747 (.Y(FE_OFN663_n4747), 
	.A(FE_OFN662_n4747));
   CLKBUFX2TS FE_OFC662_n4747 (.Y(FE_OFN662_n4747), 
	.A(FE_OFN661_n4747));
   CLKBUFX2TS FE_OFC661_n4747 (.Y(FE_OFN661_n4747), 
	.A(FE_OFN660_n4747));
   CLKBUFX2TS FE_OFC660_n4747 (.Y(FE_OFN660_n4747), 
	.A(FE_OFN659_n4747));
   CLKBUFX2TS FE_OFC659_n4747 (.Y(FE_OFN659_n4747), 
	.A(FE_OFN658_n4747));
   CLKBUFX2TS FE_OFC658_n4747 (.Y(FE_OFN658_n4747), 
	.A(FE_OFN656_n4747));
   CLKBUFX2TS FE_OFC657_n4747 (.Y(FE_OFN657_n4747), 
	.A(FE_OFN655_n4747));
   CLKBUFX2TS FE_OFC656_n4747 (.Y(FE_OFN656_n4747), 
	.A(FE_OFN654_n4747));
   CLKBUFX2TS FE_OFC655_n4747 (.Y(FE_OFN655_n4747), 
	.A(FE_OFN652_n4747));
   CLKBUFX2TS FE_OFC654_n4747 (.Y(FE_OFN654_n4747), 
	.A(FE_OFN653_n4747));
   CLKBUFX2TS FE_OFC653_n4747 (.Y(FE_OFN653_n4747), 
	.A(n4747));
   CLKBUFX2TS FE_OFC652_n4747 (.Y(FE_OFN652_n4747), 
	.A(n4747));
   CLKBUFX2TS FE_OFC651_n4741 (.Y(FE_OFN651_n4741), 
	.A(FE_OFN650_n4741));
   CLKBUFX2TS FE_OFC650_n4741 (.Y(FE_OFN650_n4741), 
	.A(FE_OFN649_n4741));
   CLKBUFX2TS FE_OFC649_n4741 (.Y(FE_OFN649_n4741), 
	.A(FE_OFN648_n4741));
   CLKBUFX2TS FE_OFC648_n4741 (.Y(FE_OFN648_n4741), 
	.A(FE_OFN647_n4741));
   CLKBUFX2TS FE_OFC647_n4741 (.Y(FE_OFN647_n4741), 
	.A(FE_OFN646_n4741));
   CLKBUFX2TS FE_OFC646_n4741 (.Y(FE_OFN646_n4741), 
	.A(FE_OFN644_n4741));
   CLKBUFX2TS FE_OFC645_n4741 (.Y(FE_OFN645_n4741), 
	.A(FE_OFN643_n4741));
   CLKBUFX2TS FE_OFC644_n4741 (.Y(FE_OFN644_n4741), 
	.A(FE_OFN640_n4741));
   CLKBUFX2TS FE_OFC643_n4741 (.Y(FE_OFN643_n4741), 
	.A(FE_OFN641_n4741));
   CLKBUFX2TS FE_OFC642_n4741 (.Y(FE_OFN642_n4741), 
	.A(FE_OFN640_n4741));
   CLKBUFX2TS FE_OFC641_n4741 (.Y(FE_OFN641_n4741), 
	.A(n4741));
   CLKBUFX2TS FE_OFC640_n4741 (.Y(FE_OFN640_n4741), 
	.A(n4741));
   CLKBUFX2TS FE_OFC639_n4742 (.Y(FE_OFN639_n4742), 
	.A(FE_OFN636_n4742));
   CLKBUFX2TS FE_OFC638_n4742 (.Y(FE_OFN638_n4742), 
	.A(FE_OFN635_n4742));
   CLKBUFX2TS FE_OFC637_n4742 (.Y(FE_OFN637_n4742), 
	.A(FE_OFN635_n4742));
   CLKBUFX2TS FE_OFC636_n4742 (.Y(FE_OFN636_n4742), 
	.A(FE_OFN633_n4742));
   CLKBUFX2TS FE_OFC635_n4742 (.Y(FE_OFN635_n4742), 
	.A(FE_OFN632_n4742));
   CLKBUFX2TS FE_OFC634_n4742 (.Y(FE_OFN634_n4742), 
	.A(FE_OFN633_n4742));
   CLKBUFX2TS FE_OFC633_n4742 (.Y(FE_OFN633_n4742), 
	.A(FE_OFN630_n4742));
   CLKBUFX2TS FE_OFC632_n4742 (.Y(FE_OFN632_n4742), 
	.A(FE_OFN631_n4742));
   CLKBUFX2TS FE_OFC631_n4742 (.Y(FE_OFN631_n4742), 
	.A(n4742));
   CLKBUFX2TS FE_OFC630_n4742 (.Y(FE_OFN630_n4742), 
	.A(n4742));
   CLKBUFX2TS FE_OFC629_n4735 (.Y(FE_OFN629_n4735), 
	.A(FE_OFN628_n4735));
   CLKBUFX2TS FE_OFC628_n4735 (.Y(FE_OFN628_n4735), 
	.A(FE_OFN627_n4735));
   CLKBUFX2TS FE_OFC627_n4735 (.Y(FE_OFN627_n4735), 
	.A(FE_OFN625_n4735));
   CLKBUFX2TS FE_OFC626_n4735 (.Y(FE_OFN626_n4735), 
	.A(FE_OFN624_n4735));
   CLKBUFX2TS FE_OFC625_n4735 (.Y(FE_OFN625_n4735), 
	.A(FE_OFN622_n4735));
   CLKBUFX2TS FE_OFC624_n4735 (.Y(FE_OFN624_n4735), 
	.A(FE_OFN623_n4735));
   CLKBUFX2TS FE_OFC623_n4735 (.Y(FE_OFN623_n4735), 
	.A(FE_OFN620_n4735));
   CLKBUFX2TS FE_OFC622_n4735 (.Y(FE_OFN622_n4735), 
	.A(FE_OFN621_n4735));
   CLKBUFX2TS FE_OFC621_n4735 (.Y(FE_OFN621_n4735), 
	.A(FE_OFN619_n4735));
   CLKBUFX2TS FE_OFC620_n4735 (.Y(FE_OFN620_n4735), 
	.A(FE_OFN619_n4735));
   CLKBUFX2TS FE_OFC619_n4735 (.Y(FE_OFN619_n4735), 
	.A(n4735));
   CLKBUFX2TS FE_OFC618_n4735 (.Y(FE_OFN618_n4735), 
	.A(n4735));
   CLKBUFX2TS FE_OFC617_n4729 (.Y(FE_OFN617_n4729), 
	.A(FE_OFN616_n4729));
   CLKBUFX2TS FE_OFC616_n4729 (.Y(FE_OFN616_n4729), 
	.A(FE_OFN615_n4729));
   CLKBUFX2TS FE_OFC615_n4729 (.Y(FE_OFN615_n4729), 
	.A(FE_OFN614_n4729));
   CLKBUFX2TS FE_OFC614_n4729 (.Y(FE_OFN614_n4729), 
	.A(FE_OFN610_n4729));
   CLKBUFX2TS FE_OFC613_n4729 (.Y(FE_OFN613_n4729), 
	.A(FE_OFN611_n4729));
   CLKBUFX2TS FE_OFC612_n4729 (.Y(FE_OFN612_n4729), 
	.A(FE_OFN611_n4729));
   CLKBUFX2TS FE_OFC611_n4729 (.Y(FE_OFN611_n4729), 
	.A(FE_OFN607_n4729));
   CLKBUFX2TS FE_OFC610_n4729 (.Y(FE_OFN610_n4729), 
	.A(FE_OFN608_n4729));
   CLKBUFX2TS FE_OFC609_n4729 (.Y(FE_OFN609_n4729), 
	.A(FE_OFN607_n4729));
   CLKBUFX2TS FE_OFC608_n4729 (.Y(FE_OFN608_n4729), 
	.A(FE_OFN606_n4729));
   CLKBUFX2TS FE_OFC607_n4729 (.Y(FE_OFN607_n4729), 
	.A(FE_OFN606_n4729));
   CLKBUFX2TS FE_OFC606_n4729 (.Y(FE_OFN606_n4729), 
	.A(n4729));
   CLKBUFX2TS FE_OFC605_n4723 (.Y(FE_OFN605_n4723), 
	.A(FE_OFN603_n4723));
   CLKBUFX2TS FE_OFC604_n4723 (.Y(FE_OFN604_n4723), 
	.A(FE_OFN603_n4723));
   CLKBUFX2TS FE_OFC603_n4723 (.Y(FE_OFN603_n4723), 
	.A(FE_OFN601_n4723));
   CLKBUFX2TS FE_OFC602_n4723 (.Y(FE_OFN602_n4723), 
	.A(FE_OFN600_n4723));
   CLKBUFX2TS FE_OFC601_n4723 (.Y(FE_OFN601_n4723), 
	.A(FE_OFN598_n4723));
   CLKBUFX2TS FE_OFC600_n4723 (.Y(FE_OFN600_n4723), 
	.A(FE_OFN597_n4723));
   CLKBUFX2TS FE_OFC599_n4723 (.Y(FE_OFN599_n4723), 
	.A(FE_OFN597_n4723));
   CLKBUFX2TS FE_OFC598_n4723 (.Y(FE_OFN598_n4723), 
	.A(FE_OFN595_n4723));
   CLKBUFX2TS FE_OFC597_n4723 (.Y(FE_OFN597_n4723), 
	.A(FE_OFN596_n4723));
   CLKBUFX2TS FE_OFC596_n4723 (.Y(FE_OFN596_n4723), 
	.A(FE_OFN594_n4723));
   CLKBUFX2TS FE_OFC595_n4723 (.Y(FE_OFN595_n4723), 
	.A(FE_OFN594_n4723));
   CLKBUFX2TS FE_OFC594_n4723 (.Y(FE_OFN594_n4723), 
	.A(n4723));
   CLKBUFX2TS FE_OFC593_n4723 (.Y(FE_OFN593_n4723), 
	.A(n4723));
   CLKBUFX2TS FE_OFC592_n4724 (.Y(FE_OFN592_n4724), 
	.A(FE_OFN591_n4724));
   CLKBUFX2TS FE_OFC591_n4724 (.Y(FE_OFN591_n4724), 
	.A(FE_OFN589_n4724));
   CLKBUFX2TS FE_OFC590_n4724 (.Y(FE_OFN590_n4724), 
	.A(FE_OFN586_n4724));
   CLKBUFX2TS FE_OFC589_n4724 (.Y(FE_OFN589_n4724), 
	.A(FE_OFN587_n4724));
   CLKBUFX2TS FE_OFC588_n4724 (.Y(FE_OFN588_n4724), 
	.A(FE_OFN586_n4724));
   CLKBUFX2TS FE_OFC587_n4724 (.Y(FE_OFN587_n4724), 
	.A(FE_OFN585_n4724));
   CLKBUFX2TS FE_OFC586_n4724 (.Y(FE_OFN586_n4724), 
	.A(FE_OFN584_n4724));
   CLKBUFX2TS FE_OFC585_n4724 (.Y(FE_OFN585_n4724), 
	.A(FE_OFN582_n4724));
   CLKBUFX2TS FE_OFC584_n4724 (.Y(FE_OFN584_n4724), 
	.A(FE_OFN583_n4724));
   CLKBUFX2TS FE_OFC583_n4724 (.Y(FE_OFN583_n4724), 
	.A(n4724));
   CLKBUFX2TS FE_OFC582_n4724 (.Y(FE_OFN582_n4724), 
	.A(n4724));
   CLKBUFX2TS FE_OFC581_n4717 (.Y(FE_OFN581_n4717), 
	.A(FE_OFN578_n4717));
   CLKBUFX2TS FE_OFC580_n4717 (.Y(FE_OFN580_n4717), 
	.A(FE_OFN578_n4717));
   CLKBUFX2TS FE_OFC579_n4717 (.Y(FE_OFN579_n4717), 
	.A(FE_OFN576_n4717));
   CLKBUFX2TS FE_OFC578_n4717 (.Y(FE_OFN578_n4717), 
	.A(FE_OFN575_n4717));
   CLKBUFX2TS FE_OFC577_n4717 (.Y(FE_OFN577_n4717), 
	.A(FE_OFN573_n4717));
   CLKBUFX2TS FE_OFC576_n4717 (.Y(FE_OFN576_n4717), 
	.A(FE_OFN574_n4717));
   CLKBUFX2TS FE_OFC575_n4717 (.Y(FE_OFN575_n4717), 
	.A(FE_OFN572_n4717));
   CLKBUFX2TS FE_OFC574_n4717 (.Y(FE_OFN574_n4717), 
	.A(FE_OFN572_n4717));
   CLKBUFX2TS FE_OFC573_n4717 (.Y(FE_OFN573_n4717), 
	.A(FE_OFN571_n4717));
   CLKBUFX2TS FE_OFC572_n4717 (.Y(FE_OFN572_n4717), 
	.A(FE_OFN570_n4717));
   CLKBUFX2TS FE_OFC571_n4717 (.Y(FE_OFN571_n4717), 
	.A(FE_OFN570_n4717));
   CLKBUFX2TS FE_OFC570_n4717 (.Y(FE_OFN570_n4717), 
	.A(n4717));
   CLKBUFX2TS FE_OFC569_n4711 (.Y(FE_OFN569_n4711), 
	.A(FE_OFN566_n4711));
   CLKBUFX2TS FE_OFC568_n4711 (.Y(FE_OFN568_n4711), 
	.A(FE_OFN564_n4711));
   CLKBUFX2TS FE_OFC567_n4711 (.Y(FE_OFN567_n4711), 
	.A(FE_OFN564_n4711));
   CLKBUFX2TS FE_OFC566_n4711 (.Y(FE_OFN566_n4711), 
	.A(FE_OFN565_n4711));
   CLKBUFX2TS FE_OFC565_n4711 (.Y(FE_OFN565_n4711), 
	.A(FE_OFN563_n4711));
   CLKBUFX2TS FE_OFC564_n4711 (.Y(FE_OFN564_n4711), 
	.A(FE_OFN561_n4711));
   CLKBUFX2TS FE_OFC563_n4711 (.Y(FE_OFN563_n4711), 
	.A(FE_OFN562_n4711));
   CLKBUFX2TS FE_OFC562_n4711 (.Y(FE_OFN562_n4711), 
	.A(FE_OFN559_n4711));
   CLKBUFX2TS FE_OFC561_n4711 (.Y(FE_OFN561_n4711), 
	.A(FE_OFN559_n4711));
   CLKBUFX2TS FE_OFC560_n4711 (.Y(FE_OFN560_n4711), 
	.A(FE_OFN559_n4711));
   CLKBUFX2TS FE_OFC559_n4711 (.Y(FE_OFN559_n4711), 
	.A(FE_OFN558_n4711));
   CLKBUFX2TS FE_OFC558_n4711 (.Y(FE_OFN558_n4711), 
	.A(n4711));
   CLKBUFX2TS FE_OFC557_n4705 (.Y(FE_OFN557_n4705), 
	.A(FE_OFN552_n4705));
   CLKBUFX2TS FE_OFC556_n4705 (.Y(FE_OFN556_n4705), 
	.A(FE_OFN551_n4705));
   CLKBUFX2TS FE_OFC555_n4705 (.Y(FE_OFN555_n4705), 
	.A(FE_OFN552_n4705));
   CLKBUFX2TS FE_OFC554_n4705 (.Y(FE_OFN554_n4705), 
	.A(FE_OFN550_n4705));
   CLKBUFX2TS FE_OFC553_n4705 (.Y(FE_OFN553_n4705), 
	.A(FE_OFN548_n4705));
   CLKBUFX2TS FE_OFC552_n4705 (.Y(FE_OFN552_n4705), 
	.A(FE_OFN548_n4705));
   CLKBUFX2TS FE_OFC551_n4705 (.Y(FE_OFN551_n4705), 
	.A(FE_OFN549_n4705));
   CLKBUFX2TS FE_OFC550_n4705 (.Y(FE_OFN550_n4705), 
	.A(FE_OFN549_n4705));
   CLKBUFX2TS FE_OFC549_n4705 (.Y(FE_OFN549_n4705), 
	.A(FE_OFN547_n4705));
   CLKBUFX2TS FE_OFC548_n4705 (.Y(FE_OFN548_n4705), 
	.A(FE_OFN547_n4705));
   CLKBUFX2TS FE_OFC547_n4705 (.Y(FE_OFN547_n4705), 
	.A(n4705));
   CLKBUFX2TS FE_OFC546_n4705 (.Y(FE_OFN546_n4705), 
	.A(n4705));
   CLKBUFX2TS FE_OFC545_n4699 (.Y(FE_OFN545_n4699), 
	.A(FE_OFN541_n4699));
   CLKBUFX2TS FE_OFC544_n4699 (.Y(FE_OFN544_n4699), 
	.A(FE_OFN542_n4699));
   CLKBUFX2TS FE_OFC543_n4699 (.Y(FE_OFN543_n4699), 
	.A(FE_OFN541_n4699));
   CLKBUFX2TS FE_OFC542_n4699 (.Y(FE_OFN542_n4699), 
	.A(FE_OFN539_n4699));
   CLKBUFX2TS FE_OFC541_n4699 (.Y(FE_OFN541_n4699), 
	.A(FE_OFN540_n4699));
   CLKBUFX2TS FE_OFC540_n4699 (.Y(FE_OFN540_n4699), 
	.A(FE_OFN537_n4699));
   CLKBUFX2TS FE_OFC539_n4699 (.Y(FE_OFN539_n4699), 
	.A(FE_OFN536_n4699));
   CLKBUFX2TS FE_OFC538_n4699 (.Y(FE_OFN538_n4699), 
	.A(FE_OFN536_n4699));
   CLKBUFX2TS FE_OFC537_n4699 (.Y(FE_OFN537_n4699), 
	.A(FE_OFN535_n4699));
   CLKBUFX2TS FE_OFC536_n4699 (.Y(FE_OFN536_n4699), 
	.A(FE_OFN535_n4699));
   CLKBUFX2TS FE_OFC535_n4699 (.Y(FE_OFN535_n4699), 
	.A(n4699));
   CLKBUFX2TS FE_OFC534_n4699 (.Y(FE_OFN534_n4699), 
	.A(n4699));
   CLKBUFX2TS FE_OFC533_n4700 (.Y(FE_OFN533_n4700), 
	.A(FE_OFN531_n4700));
   CLKBUFX2TS FE_OFC532_n4700 (.Y(FE_OFN532_n4700), 
	.A(FE_OFN530_n4700));
   CLKBUFX2TS FE_OFC531_n4700 (.Y(FE_OFN531_n4700), 
	.A(FE_OFN529_n4700));
   CLKBUFX2TS FE_OFC530_n4700 (.Y(FE_OFN530_n4700), 
	.A(FE_OFN528_n4700));
   CLKBUFX2TS FE_OFC529_n4700 (.Y(FE_OFN529_n4700), 
	.A(FE_OFN526_n4700));
   CLKBUFX2TS FE_OFC528_n4700 (.Y(FE_OFN528_n4700), 
	.A(FE_OFN527_n4700));
   CLKBUFX2TS FE_OFC527_n4700 (.Y(FE_OFN527_n4700), 
	.A(FE_OFN525_n4700));
   CLKBUFX2TS FE_OFC526_n4700 (.Y(FE_OFN526_n4700), 
	.A(FE_OFN524_n4700));
   CLKBUFX2TS FE_OFC525_n4700 (.Y(FE_OFN525_n4700), 
	.A(FE_OFN523_n4700));
   CLKBUFX2TS FE_OFC524_n4700 (.Y(FE_OFN524_n4700), 
	.A(FE_OFN523_n4700));
   CLKBUFX2TS FE_OFC523_n4700 (.Y(FE_OFN523_n4700), 
	.A(n4700));
   CLKBUFX2TS FE_OFC522_n4693 (.Y(FE_OFN522_n4693), 
	.A(FE_OFN521_n4693));
   CLKBUFX2TS FE_OFC521_n4693 (.Y(FE_OFN521_n4693), 
	.A(FE_OFN520_n4693));
   CLKBUFX2TS FE_OFC520_n4693 (.Y(FE_OFN520_n4693), 
	.A(FE_OFN519_n4693));
   CLKBUFX2TS FE_OFC519_n4693 (.Y(FE_OFN519_n4693), 
	.A(FE_OFN518_n4693));
   CLKBUFX2TS FE_OFC518_n4693 (.Y(FE_OFN518_n4693), 
	.A(FE_OFN517_n4693));
   CLKBUFX2TS FE_OFC517_n4693 (.Y(FE_OFN517_n4693), 
	.A(FE_OFN516_n4693));
   CLKBUFX2TS FE_OFC516_n4693 (.Y(FE_OFN516_n4693), 
	.A(FE_OFN515_n4693));
   CLKBUFX2TS FE_OFC515_n4693 (.Y(FE_OFN515_n4693), 
	.A(FE_OFN513_n4693));
   CLKBUFX2TS FE_OFC514_n4693 (.Y(FE_OFN514_n4693), 
	.A(FE_OFN513_n4693));
   CLKBUFX2TS FE_OFC513_n4693 (.Y(FE_OFN513_n4693), 
	.A(FE_OFN512_n4693));
   CLKBUFX2TS FE_OFC512_n4693 (.Y(FE_OFN512_n4693), 
	.A(FE_OFN511_n4693));
   CLKBUFX2TS FE_OFC511_n4693 (.Y(FE_OFN511_n4693), 
	.A(n4693));
   CLKBUFX2TS FE_OFC510_n8055 (.Y(FE_OFN510_n8055), 
	.A(FE_OFN509_n8055));
   CLKBUFX2TS FE_OFC509_n8055 (.Y(FE_OFN509_n8055), 
	.A(FE_OFN508_n8055));
   CLKBUFX2TS FE_OFC508_n8055 (.Y(FE_OFN508_n8055), 
	.A(n8055));
   CLKBUFX2TS FE_OFC507_n4681 (.Y(FE_OFN507_n4681), 
	.A(FE_OFN505_n4681));
   CLKBUFX2TS FE_OFC506_n4681 (.Y(FE_OFN506_n4681), 
	.A(FE_OFN504_n4681));
   CLKBUFX2TS FE_OFC505_n4681 (.Y(FE_OFN505_n4681), 
	.A(FE_OFN503_n4681));
   CLKBUFX2TS FE_OFC504_n4681 (.Y(FE_OFN504_n4681), 
	.A(FE_OFN503_n4681));
   CLKBUFX2TS FE_OFC503_n4681 (.Y(FE_OFN503_n4681), 
	.A(FE_OFN502_n4681));
   CLKBUFX2TS FE_OFC502_n4681 (.Y(FE_OFN502_n4681), 
	.A(FE_OFN501_n4681));
   CLKBUFX2TS FE_OFC501_n4681 (.Y(FE_OFN501_n4681), 
	.A(FE_OFN500_n4681));
   CLKBUFX2TS FE_OFC500_n4681 (.Y(FE_OFN500_n4681), 
	.A(FE_OFN499_n4681));
   CLKBUFX2TS FE_OFC499_n4681 (.Y(FE_OFN499_n4681), 
	.A(FE_OFN498_n4681));
   CLKBUFX2TS FE_OFC498_n4681 (.Y(FE_OFN498_n4681), 
	.A(FE_OFN497_n4681));
   CLKBUFX2TS FE_OFC497_n4681 (.Y(FE_OFN497_n4681), 
	.A(n4681));
   CLKBUFX2TS FE_OFC496_n4681 (.Y(FE_OFN496_n4681), 
	.A(n4681));
   CLKBUFX2TS FE_OFC495_n4682 (.Y(FE_OFN495_n4682), 
	.A(FE_OFN491_n4682));
   CLKBUFX2TS FE_OFC494_n4682 (.Y(FE_OFN494_n4682), 
	.A(FE_OFN492_n4682));
   CLKBUFX2TS FE_OFC493_n4682 (.Y(FE_OFN493_n4682), 
	.A(FE_OFN492_n4682));
   CLKBUFX2TS FE_OFC492_n4682 (.Y(FE_OFN492_n4682), 
	.A(FE_OFN490_n4682));
   CLKBUFX2TS FE_OFC491_n4682 (.Y(FE_OFN491_n4682), 
	.A(FE_OFN487_n4682));
   CLKBUFX2TS FE_OFC490_n4682 (.Y(FE_OFN490_n4682), 
	.A(FE_OFN488_n4682));
   CLKBUFX2TS FE_OFC489_n4682 (.Y(FE_OFN489_n4682), 
	.A(FE_OFN486_n4682));
   CLKBUFX2TS FE_OFC488_n4682 (.Y(FE_OFN488_n4682), 
	.A(n4682));
   CLKBUFX2TS FE_OFC487_n4682 (.Y(FE_OFN487_n4682), 
	.A(FE_OFN486_n4682));
   CLKBUFX2TS FE_OFC486_n4682 (.Y(FE_OFN486_n4682), 
	.A(n4682));
   CLKBUFX2TS FE_OFC485_n4675 (.Y(FE_OFN485_n4675), 
	.A(FE_OFN483_n4675));
   CLKBUFX2TS FE_OFC484_n4675 (.Y(FE_OFN484_n4675), 
	.A(FE_OFN483_n4675));
   CLKBUFX2TS FE_OFC483_n4675 (.Y(FE_OFN483_n4675), 
	.A(FE_OFN482_n4675));
   CLKBUFX2TS FE_OFC482_n4675 (.Y(FE_OFN482_n4675), 
	.A(FE_OFN481_n4675));
   CLKBUFX2TS FE_OFC481_n4675 (.Y(FE_OFN481_n4675), 
	.A(FE_OFN479_n4675));
   CLKBUFX2TS FE_OFC480_n4675 (.Y(FE_OFN480_n4675), 
	.A(FE_OFN479_n4675));
   CLKBUFX2TS FE_OFC479_n4675 (.Y(FE_OFN479_n4675), 
	.A(FE_OFN478_n4675));
   CLKBUFX2TS FE_OFC478_n4675 (.Y(FE_OFN478_n4675), 
	.A(FE_OFN477_n4675));
   CLKBUFX2TS FE_OFC477_n4675 (.Y(FE_OFN477_n4675), 
	.A(FE_OFN476_n4675));
   CLKBUFX2TS FE_OFC476_n4675 (.Y(FE_OFN476_n4675), 
	.A(FE_OFN475_n4675));
   CLKBUFX2TS FE_OFC475_n4675 (.Y(FE_OFN475_n4675), 
	.A(FE_OFN474_n4675));
   CLKBUFX2TS FE_OFC474_n4675 (.Y(FE_OFN474_n4675), 
	.A(n4675));
   CLKBUFX2TS FE_OFC473_n4676 (.Y(FE_OFN473_n4676), 
	.A(FE_OFN471_n4676));
   CLKBUFX2TS FE_OFC472_n4676 (.Y(FE_OFN472_n4676), 
	.A(FE_OFN471_n4676));
   CLKBUFX2TS FE_OFC471_n4676 (.Y(FE_OFN471_n4676), 
	.A(FE_OFN468_n4676));
   CLKBUFX2TS FE_OFC470_n4676 (.Y(FE_OFN470_n4676), 
	.A(FE_OFN467_n4676));
   CLKBUFX2TS FE_OFC469_n4676 (.Y(FE_OFN469_n4676), 
	.A(FE_OFN467_n4676));
   CLKBUFX2TS FE_OFC468_n4676 (.Y(FE_OFN468_n4676), 
	.A(FE_OFN466_n4676));
   CLKBUFX2TS FE_OFC467_n4676 (.Y(FE_OFN467_n4676), 
	.A(FE_OFN465_n4676));
   CLKBUFX2TS FE_OFC466_n4676 (.Y(FE_OFN466_n4676), 
	.A(FE_OFN464_n4676));
   CLKBUFX2TS FE_OFC465_n4676 (.Y(FE_OFN465_n4676), 
	.A(FE_OFN463_n4676));
   CLKBUFX2TS FE_OFC464_n4676 (.Y(FE_OFN464_n4676), 
	.A(FE_OFN463_n4676));
   CLKBUFX2TS FE_OFC463_n4676 (.Y(FE_OFN463_n4676), 
	.A(n4676));
   CLKBUFX2TS FE_OFC462_n4688 (.Y(FE_OFN462_n4688), 
	.A(FE_OFN460_n4688));
   CLKBUFX2TS FE_OFC461_n4688 (.Y(FE_OFN461_n4688), 
	.A(FE_OFN459_n4688));
   CLKBUFX2TS FE_OFC460_n4688 (.Y(FE_OFN460_n4688), 
	.A(FE_OFN459_n4688));
   CLKBUFX2TS FE_OFC459_n4688 (.Y(FE_OFN459_n4688), 
	.A(FE_OFN458_n4688));
   CLKBUFX2TS FE_OFC458_n4688 (.Y(FE_OFN458_n4688), 
	.A(FE_OFN457_n4688));
   CLKBUFX2TS FE_OFC457_n4688 (.Y(FE_OFN457_n4688), 
	.A(FE_OFN456_n4688));
   CLKBUFX2TS FE_OFC456_n4688 (.Y(FE_OFN456_n4688), 
	.A(FE_OFN454_n4688));
   CLKBUFX2TS FE_OFC455_n4688 (.Y(FE_OFN455_n4688), 
	.A(FE_OFN453_n4688));
   CLKBUFX2TS FE_OFC454_n4688 (.Y(FE_OFN454_n4688), 
	.A(n4688));
   CLKBUFX2TS FE_OFC453_n4688 (.Y(FE_OFN453_n4688), 
	.A(n4688));
   CLKBUFX2TS FE_OFC452_n4694 (.Y(FE_OFN452_n4694), 
	.A(FE_OFN450_n4694));
   CLKBUFX2TS FE_OFC451_n4694 (.Y(FE_OFN451_n4694), 
	.A(FE_OFN450_n4694));
   CLKBUFX2TS FE_OFC450_n4694 (.Y(FE_OFN450_n4694), 
	.A(FE_OFN448_n4694));
   CLKBUFX2TS FE_OFC449_n4694 (.Y(FE_OFN449_n4694), 
	.A(FE_OFN447_n4694));
   CLKBUFX2TS FE_OFC448_n4694 (.Y(FE_OFN448_n4694), 
	.A(FE_OFN445_n4694));
   CLKBUFX2TS FE_OFC447_n4694 (.Y(FE_OFN447_n4694), 
	.A(FE_OFN446_n4694));
   CLKBUFX2TS FE_OFC446_n4694 (.Y(FE_OFN446_n4694), 
	.A(FE_OFN444_n4694));
   CLKBUFX2TS FE_OFC445_n4694 (.Y(FE_OFN445_n4694), 
	.A(FE_OFN443_n4694));
   CLKBUFX2TS FE_OFC444_n4694 (.Y(FE_OFN444_n4694), 
	.A(n4694));
   CLKBUFX2TS FE_OFC443_n4694 (.Y(FE_OFN443_n4694), 
	.A(n4694));
   CLKBUFX2TS FE_OFC442_n4706 (.Y(FE_OFN442_n4706), 
	.A(FE_OFN438_n4706));
   CLKBUFX2TS FE_OFC441_n4706 (.Y(FE_OFN441_n4706), 
	.A(FE_OFN438_n4706));
   CLKBUFX2TS FE_OFC440_n4706 (.Y(FE_OFN440_n4706), 
	.A(FE_OFN435_n4706));
   CLKBUFX2TS FE_OFC439_n4706 (.Y(FE_OFN439_n4706), 
	.A(FE_OFN436_n4706));
   CLKBUFX2TS FE_OFC438_n4706 (.Y(FE_OFN438_n4706), 
	.A(FE_OFN434_n4706));
   CLKBUFX2TS FE_OFC437_n4706 (.Y(FE_OFN437_n4706), 
	.A(FE_OFN434_n4706));
   CLKBUFX2TS FE_OFC436_n4706 (.Y(FE_OFN436_n4706), 
	.A(FE_OFN433_n4706));
   CLKBUFX2TS FE_OFC435_n4706 (.Y(FE_OFN435_n4706), 
	.A(FE_OFN433_n4706));
   CLKBUFX2TS FE_OFC434_n4706 (.Y(FE_OFN434_n4706), 
	.A(n4706));
   CLKBUFX2TS FE_OFC433_n4706 (.Y(FE_OFN433_n4706), 
	.A(n4706));
   CLKBUFX2TS FE_OFC432_n4712 (.Y(FE_OFN432_n4712), 
	.A(FE_OFN429_n4712));
   CLKBUFX2TS FE_OFC431_n4712 (.Y(FE_OFN431_n4712), 
	.A(FE_OFN427_n4712));
   CLKBUFX2TS FE_OFC430_n4712 (.Y(FE_OFN430_n4712), 
	.A(FE_OFN427_n4712));
   CLKBUFX2TS FE_OFC429_n4712 (.Y(FE_OFN429_n4712), 
	.A(FE_OFN428_n4712));
   CLKBUFX2TS FE_OFC428_n4712 (.Y(FE_OFN428_n4712), 
	.A(FE_OFN426_n4712));
   CLKBUFX2TS FE_OFC427_n4712 (.Y(FE_OFN427_n4712), 
	.A(FE_OFN425_n4712));
   CLKBUFX2TS FE_OFC426_n4712 (.Y(FE_OFN426_n4712), 
	.A(FE_OFN424_n4712));
   CLKBUFX2TS FE_OFC425_n4712 (.Y(FE_OFN425_n4712), 
	.A(FE_OFN424_n4712));
   CLKBUFX2TS FE_OFC424_n4712 (.Y(FE_OFN424_n4712), 
	.A(FE_OFN423_n4712));
   CLKBUFX2TS FE_OFC423_n4712 (.Y(FE_OFN423_n4712), 
	.A(n4712));
   CLKBUFX2TS FE_OFC422_n3776 (.Y(FE_OFN422_n3776), 
	.A(FE_OFN420_n3776));
   CLKBUFX2TS FE_OFC421_n3776 (.Y(FE_OFN421_n3776), 
	.A(FE_OFN420_n3776));
   CLKBUFX2TS FE_OFC420_n3776 (.Y(FE_OFN420_n3776), 
	.A(FE_OFN418_n3776));
   CLKBUFX2TS FE_OFC419_n3776 (.Y(FE_OFN419_n3776), 
	.A(FE_OFN417_n3776));
   CLKBUFX2TS FE_OFC418_n3776 (.Y(FE_OFN418_n3776), 
	.A(FE_OFN416_n3776));
   CLKBUFX2TS FE_OFC417_n3776 (.Y(FE_OFN417_n3776), 
	.A(FE_OFN416_n3776));
   CLKBUFX2TS FE_OFC416_n3776 (.Y(FE_OFN416_n3776), 
	.A(FE_OFN415_n3776));
   CLKBUFX2TS FE_OFC415_n3776 (.Y(FE_OFN415_n3776), 
	.A(FE_OFN413_n3776));
   CLKBUFX2TS FE_OFC414_n3776 (.Y(FE_OFN414_n3776), 
	.A(FE_OFN413_n3776));
   CLKBUFX2TS FE_OFC413_n3776 (.Y(FE_OFN413_n3776), 
	.A(FE_OFN412_n3776));
   CLKBUFX2TS FE_OFC412_n3776 (.Y(FE_OFN412_n3776), 
	.A(n3776));
   CLKBUFX2TS FE_OFC411_n3777 (.Y(FE_OFN411_n3777), 
	.A(FE_OFN409_n3777));
   CLKBUFX2TS FE_OFC410_n3777 (.Y(FE_OFN410_n3777), 
	.A(FE_OFN407_n3777));
   CLKBUFX2TS FE_OFC409_n3777 (.Y(FE_OFN409_n3777), 
	.A(FE_OFN406_n3777));
   CLKBUFX2TS FE_OFC408_n3777 (.Y(FE_OFN408_n3777), 
	.A(FE_OFN407_n3777));
   CLKBUFX2TS FE_OFC407_n3777 (.Y(FE_OFN407_n3777), 
	.A(FE_OFN404_n3777));
   CLKBUFX2TS FE_OFC406_n3777 (.Y(FE_OFN406_n3777), 
	.A(FE_OFN403_n3777));
   CLKBUFX2TS FE_OFC405_n3777 (.Y(FE_OFN405_n3777), 
	.A(FE_OFN401_n3777));
   CLKBUFX2TS FE_OFC404_n3777 (.Y(FE_OFN404_n3777), 
	.A(FE_OFN402_n3777));
   CLKBUFX2TS FE_OFC403_n3777 (.Y(FE_OFN403_n3777), 
	.A(FE_OFN402_n3777));
   CLKBUFX2TS FE_OFC402_n3777 (.Y(FE_OFN402_n3777), 
	.A(n3777));
   CLKBUFX2TS FE_OFC401_n3777 (.Y(FE_OFN401_n3777), 
	.A(n3777));
   CLKBUFX2TS FE_OFC400_n4718 (.Y(FE_OFN400_n4718), 
	.A(FE_OFN396_n4718));
   CLKBUFX2TS FE_OFC399_n4718 (.Y(FE_OFN399_n4718), 
	.A(FE_OFN395_n4718));
   CLKBUFX2TS FE_OFC398_n4718 (.Y(FE_OFN398_n4718), 
	.A(FE_OFN395_n4718));
   CLKBUFX2TS FE_OFC397_n4718 (.Y(FE_OFN397_n4718), 
	.A(FE_OFN394_n4718));
   CLKBUFX2TS FE_OFC396_n4718 (.Y(FE_OFN396_n4718), 
	.A(FE_OFN394_n4718));
   CLKBUFX2TS FE_OFC395_n4718 (.Y(FE_OFN395_n4718), 
	.A(FE_OFN392_n4718));
   CLKBUFX2TS FE_OFC394_n4718 (.Y(FE_OFN394_n4718), 
	.A(FE_OFN393_n4718));
   CLKBUFX2TS FE_OFC393_n4718 (.Y(FE_OFN393_n4718), 
	.A(FE_OFN390_n4718));
   CLKBUFX2TS FE_OFC392_n4718 (.Y(FE_OFN392_n4718), 
	.A(FE_OFN390_n4718));
   CLKBUFX2TS FE_OFC391_n4718 (.Y(FE_OFN391_n4718), 
	.A(FE_OFN390_n4718));
   CLKBUFX2TS FE_OFC390_n4718 (.Y(FE_OFN390_n4718), 
	.A(n4718));
   CLKBUFX2TS FE_OFC389_n4730 (.Y(FE_OFN389_n4730), 
	.A(FE_OFN387_n4730));
   CLKBUFX2TS FE_OFC388_n4730 (.Y(FE_OFN388_n4730), 
	.A(FE_OFN386_n4730));
   CLKBUFX2TS FE_OFC387_n4730 (.Y(FE_OFN387_n4730), 
	.A(FE_OFN384_n4730));
   CLKBUFX2TS FE_OFC386_n4730 (.Y(FE_OFN386_n4730), 
	.A(FE_OFN385_n4730));
   CLKBUFX2TS FE_OFC385_n4730 (.Y(FE_OFN385_n4730), 
	.A(FE_OFN382_n4730));
   CLKBUFX2TS FE_OFC384_n4730 (.Y(FE_OFN384_n4730), 
	.A(FE_OFN383_n4730));
   CLKBUFX2TS FE_OFC383_n4730 (.Y(FE_OFN383_n4730), 
	.A(FE_OFN381_n4730));
   CLKBUFX2TS FE_OFC382_n4730 (.Y(FE_OFN382_n4730), 
	.A(FE_OFN380_n4730));
   CLKBUFX2TS FE_OFC381_n4730 (.Y(FE_OFN381_n4730), 
	.A(FE_OFN379_n4730));
   CLKBUFX2TS FE_OFC380_n4730 (.Y(FE_OFN380_n4730), 
	.A(FE_OFN379_n4730));
   CLKBUFX2TS FE_OFC379_n4730 (.Y(FE_OFN379_n4730), 
	.A(n4730));
   CLKBUFX2TS FE_OFC378_n4736 (.Y(FE_OFN378_n4736), 
	.A(FE_OFN376_n4736));
   CLKBUFX2TS FE_OFC377_n4736 (.Y(FE_OFN377_n4736), 
	.A(FE_OFN375_n4736));
   CLKBUFX2TS FE_OFC376_n4736 (.Y(FE_OFN376_n4736), 
	.A(FE_OFN374_n4736));
   CLKBUFX2TS FE_OFC375_n4736 (.Y(FE_OFN375_n4736), 
	.A(FE_OFN373_n4736));
   CLKBUFX2TS FE_OFC374_n4736 (.Y(FE_OFN374_n4736), 
	.A(FE_OFN371_n4736));
   CLKBUFX2TS FE_OFC373_n4736 (.Y(FE_OFN373_n4736), 
	.A(FE_OFN372_n4736));
   CLKBUFX2TS FE_OFC372_n4736 (.Y(FE_OFN372_n4736), 
	.A(FE_OFN370_n4736));
   CLKBUFX2TS FE_OFC371_n4736 (.Y(FE_OFN371_n4736), 
	.A(FE_OFN369_n4736));
   CLKBUFX2TS FE_OFC370_n4736 (.Y(FE_OFN370_n4736), 
	.A(n4736));
   CLKBUFX2TS FE_OFC369_n4736 (.Y(FE_OFN369_n4736), 
	.A(n4736));
   CLKBUFX2TS FE_OFC368_n4748 (.Y(FE_OFN368_n4748), 
	.A(FE_OFN366_n4748));
   CLKBUFX2TS FE_OFC367_n4748 (.Y(FE_OFN367_n4748), 
	.A(FE_OFN364_n4748));
   CLKBUFX2TS FE_OFC366_n4748 (.Y(FE_OFN366_n4748), 
	.A(FE_OFN363_n4748));
   CLKBUFX2TS FE_OFC365_n4748 (.Y(FE_OFN365_n4748), 
	.A(FE_OFN364_n4748));
   CLKBUFX2TS FE_OFC364_n4748 (.Y(FE_OFN364_n4748), 
	.A(FE_OFN362_n4748));
   CLKBUFX2TS FE_OFC363_n4748 (.Y(FE_OFN363_n4748), 
	.A(FE_OFN361_n4748));
   CLKBUFX2TS FE_OFC362_n4748 (.Y(FE_OFN362_n4748), 
	.A(FE_OFN359_n4748));
   CLKBUFX2TS FE_OFC361_n4748 (.Y(FE_OFN361_n4748), 
	.A(FE_OFN360_n4748));
   CLKBUFX2TS FE_OFC360_n4748 (.Y(FE_OFN360_n4748), 
	.A(n4748));
   CLKBUFX2TS FE_OFC359_n4748 (.Y(FE_OFN359_n4748), 
	.A(n4748));
   CLKBUFX2TS FE_OFC358_n4754 (.Y(FE_OFN358_n4754), 
	.A(FE_OFN357_n4754));
   CLKBUFX2TS FE_OFC357_n4754 (.Y(FE_OFN357_n4754), 
	.A(FE_OFN356_n4754));
   CLKBUFX2TS FE_OFC356_n4754 (.Y(FE_OFN356_n4754), 
	.A(FE_OFN355_n4754));
   CLKBUFX2TS FE_OFC355_n4754 (.Y(FE_OFN355_n4754), 
	.A(FE_OFN354_n4754));
   CLKBUFX2TS FE_OFC354_n4754 (.Y(FE_OFN354_n4754), 
	.A(FE_OFN352_n4754));
   CLKBUFX2TS FE_OFC353_n4754 (.Y(FE_OFN353_n4754), 
	.A(FE_OFN350_n4754));
   CLKBUFX2TS FE_OFC352_n4754 (.Y(FE_OFN352_n4754), 
	.A(FE_OFN351_n4754));
   CLKBUFX2TS FE_OFC351_n4754 (.Y(FE_OFN351_n4754), 
	.A(FE_OFN349_n4754));
   CLKBUFX2TS FE_OFC350_n4754 (.Y(FE_OFN350_n4754), 
	.A(n4754));
   CLKBUFX2TS FE_OFC349_n4754 (.Y(FE_OFN349_n4754), 
	.A(n4754));
   CLKBUFX2TS FE_OFC348_n4760 (.Y(FE_OFN348_n4760), 
	.A(FE_OFN345_n4760));
   CLKBUFX2TS FE_OFC347_n4760 (.Y(FE_OFN347_n4760), 
	.A(FE_OFN345_n4760));
   CLKBUFX2TS FE_OFC346_n4760 (.Y(FE_OFN346_n4760), 
	.A(FE_OFN343_n4760));
   CLKBUFX2TS FE_OFC345_n4760 (.Y(FE_OFN345_n4760), 
	.A(FE_OFN342_n4760));
   CLKBUFX2TS FE_OFC344_n4760 (.Y(FE_OFN344_n4760), 
	.A(FE_OFN343_n4760));
   CLKBUFX2TS FE_OFC343_n4760 (.Y(FE_OFN343_n4760), 
	.A(FE_OFN339_n4760));
   CLKBUFX2TS FE_OFC342_n4760 (.Y(FE_OFN342_n4760), 
	.A(FE_OFN338_n4760));
   CLKBUFX2TS FE_OFC341_n4760 (.Y(FE_OFN341_n4760), 
	.A(FE_OFN339_n4760));
   CLKBUFX2TS FE_OFC340_n4760 (.Y(FE_OFN340_n4760), 
	.A(FE_OFN338_n4760));
   CLKBUFX2TS FE_OFC339_n4760 (.Y(FE_OFN339_n4760), 
	.A(n4760));
   CLKBUFX2TS FE_OFC338_n4760 (.Y(FE_OFN338_n4760), 
	.A(n4760));
   CLKBUFX2TS FE_OFC337_n4573 (.Y(FE_OFN337_n4573), 
	.A(FE_OFN336_n4573));
   CLKBUFX2TS FE_OFC336_n4573 (.Y(FE_OFN336_n4573), 
	.A(FE_OFN335_n4573));
   CLKBUFX2TS FE_OFC335_n4573 (.Y(FE_OFN335_n4573), 
	.A(FE_OFN334_n4573));
   CLKBUFX2TS FE_OFC334_n4573 (.Y(FE_OFN334_n4573), 
	.A(FE_OFN333_n4573));
   CLKBUFX2TS FE_OFC333_n4573 (.Y(FE_OFN333_n4573), 
	.A(FE_OFN332_n4573));
   CLKBUFX2TS FE_OFC332_n4573 (.Y(FE_OFN332_n4573), 
	.A(FE_OFN331_n4573));
   CLKBUFX2TS FE_OFC331_n4573 (.Y(FE_OFN331_n4573), 
	.A(FE_OFN329_n4573));
   CLKBUFX2TS FE_OFC330_n4573 (.Y(FE_OFN330_n4573), 
	.A(FE_OFN329_n4573));
   CLKBUFX2TS FE_OFC329_n4573 (.Y(FE_OFN329_n4573), 
	.A(FE_OFN328_n4573));
   CLKBUFX2TS FE_OFC328_n4573 (.Y(FE_OFN328_n4573), 
	.A(FE_OFN327_n4573));
   CLKBUFX2TS FE_OFC327_n4573 (.Y(FE_OFN327_n4573), 
	.A(n4573));
   CLKBUFX2TS FE_OFC326_n8056 (.Y(FE_OFN326_n8056), 
	.A(FE_OFN325_n8056));
   CLKBUFX2TS FE_OFC325_n8056 (.Y(FE_OFN325_n8056), 
	.A(n8056));
   CLKBUFX2TS FE_OFC324_n4561 (.Y(FE_OFN324_n4561), 
	.A(FE_OFN323_n4561));
   CLKBUFX2TS FE_OFC323_n4561 (.Y(FE_OFN323_n4561), 
	.A(FE_OFN322_n4561));
   CLKBUFX2TS FE_OFC322_n4561 (.Y(FE_OFN322_n4561), 
	.A(FE_OFN319_n4561));
   CLKBUFX2TS FE_OFC321_n4561 (.Y(FE_OFN321_n4561), 
	.A(FE_OFN318_n4561));
   CLKBUFX2TS FE_OFC320_n4561 (.Y(FE_OFN320_n4561), 
	.A(FE_OFN315_n4561));
   CLKBUFX2TS FE_OFC319_n4561 (.Y(FE_OFN319_n4561), 
	.A(FE_OFN317_n4561));
   CLKBUFX2TS FE_OFC318_n4561 (.Y(FE_OFN318_n4561), 
	.A(FE_OFN317_n4561));
   CLKBUFX2TS FE_OFC317_n4561 (.Y(FE_OFN317_n4561), 
	.A(FE_OFN316_n4561));
   CLKBUFX2TS FE_OFC316_n4561 (.Y(FE_OFN316_n4561), 
	.A(FE_OFN314_n4561));
   CLKBUFX2TS FE_OFC315_n4561 (.Y(FE_OFN315_n4561), 
	.A(FE_OFN314_n4561));
   CLKBUFX2TS FE_OFC314_n4561 (.Y(FE_OFN314_n4561), 
	.A(FE_OFN313_n4561));
   CLKBUFX2TS FE_OFC313_n4561 (.Y(FE_OFN313_n4561), 
	.A(n4561));
   CLKBUFX2TS FE_OFC312_n4555 (.Y(FE_OFN312_n4555), 
	.A(FE_OFN311_n4555));
   CLKBUFX2TS FE_OFC311_n4555 (.Y(FE_OFN311_n4555), 
	.A(FE_OFN310_n4555));
   CLKBUFX2TS FE_OFC310_n4555 (.Y(FE_OFN310_n4555), 
	.A(FE_OFN306_n4555));
   CLKBUFX2TS FE_OFC309_n4555 (.Y(FE_OFN309_n4555), 
	.A(FE_OFN307_n4555));
   CLKBUFX2TS FE_OFC308_n4555 (.Y(FE_OFN308_n4555), 
	.A(FE_OFN305_n4555));
   CLKBUFX2TS FE_OFC307_n4555 (.Y(FE_OFN307_n4555), 
	.A(FE_OFN305_n4555));
   CLKBUFX2TS FE_OFC306_n4555 (.Y(FE_OFN306_n4555), 
	.A(FE_OFN304_n4555));
   CLKBUFX2TS FE_OFC305_n4555 (.Y(FE_OFN305_n4555), 
	.A(FE_OFN303_n4555));
   CLKBUFX2TS FE_OFC304_n4555 (.Y(FE_OFN304_n4555), 
	.A(FE_OFN303_n4555));
   CLKBUFX2TS FE_OFC303_n4555 (.Y(FE_OFN303_n4555), 
	.A(FE_OFN302_n4555));
   CLKBUFX2TS FE_OFC302_n4555 (.Y(FE_OFN302_n4555), 
	.A(FE_OFN301_n4555));
   CLKBUFX2TS FE_OFC301_n4555 (.Y(FE_OFN301_n4555), 
	.A(n4555));
   CLKBUFX2TS FE_OFC300_n4556 (.Y(FE_OFN300_n4556), 
	.A(FE_OFN298_n4556));
   CLKBUFX2TS FE_OFC299_n4556 (.Y(FE_OFN299_n4556), 
	.A(FE_OFN294_n4556));
   CLKBUFX2TS FE_OFC298_n4556 (.Y(FE_OFN298_n4556), 
	.A(FE_OFN294_n4556));
   CLKBUFX2TS FE_OFC297_n4556 (.Y(FE_OFN297_n4556), 
	.A(FE_OFN293_n4556));
   CLKBUFX2TS FE_OFC296_n4556 (.Y(FE_OFN296_n4556), 
	.A(FE_OFN293_n4556));
   CLKBUFX2TS FE_OFC295_n4556 (.Y(FE_OFN295_n4556), 
	.A(FE_OFN292_n4556));
   CLKBUFX2TS FE_OFC294_n4556 (.Y(FE_OFN294_n4556), 
	.A(FE_OFN291_n4556));
   CLKBUFX2TS FE_OFC293_n4556 (.Y(FE_OFN293_n4556), 
	.A(FE_OFN292_n4556));
   CLKBUFX2TS FE_OFC292_n4556 (.Y(FE_OFN292_n4556), 
	.A(FE_OFN291_n4556));
   CLKBUFX2TS FE_OFC291_n4556 (.Y(FE_OFN291_n4556), 
	.A(n4556));
   CLKBUFX2TS FE_OFC290_n4549 (.Y(FE_OFN290_n4549), 
	.A(FE_OFN289_n4549));
   CLKBUFX2TS FE_OFC289_n4549 (.Y(FE_OFN289_n4549), 
	.A(FE_OFN288_n4549));
   CLKBUFX2TS FE_OFC288_n4549 (.Y(FE_OFN288_n4549), 
	.A(FE_OFN287_n4549));
   CLKBUFX2TS FE_OFC287_n4549 (.Y(FE_OFN287_n4549), 
	.A(FE_OFN286_n4549));
   CLKBUFX2TS FE_OFC286_n4549 (.Y(FE_OFN286_n4549), 
	.A(FE_OFN285_n4549));
   CLKBUFX2TS FE_OFC285_n4549 (.Y(FE_OFN285_n4549), 
	.A(FE_OFN284_n4549));
   CLKBUFX2TS FE_OFC284_n4549 (.Y(FE_OFN284_n4549), 
	.A(FE_OFN283_n4549));
   CLKBUFX2TS FE_OFC283_n4549 (.Y(FE_OFN283_n4549), 
	.A(FE_OFN282_n4549));
   CLKBUFX2TS FE_OFC282_n4549 (.Y(FE_OFN282_n4549), 
	.A(FE_OFN280_n4549));
   CLKBUFX2TS FE_OFC281_n4549 (.Y(FE_OFN281_n4549), 
	.A(FE_OFN279_n4549));
   CLKBUFX2TS FE_OFC280_n4549 (.Y(FE_OFN280_n4549), 
	.A(FE_OFN279_n4549));
   CLKBUFX2TS FE_OFC279_n4549 (.Y(FE_OFN279_n4549), 
	.A(n4549));
   CLKBUFX2TS FE_OFC278_n4543 (.Y(FE_OFN278_n4543), 
	.A(FE_OFN276_n4543));
   CLKBUFX2TS FE_OFC277_n4543 (.Y(FE_OFN277_n4543), 
	.A(FE_OFN275_n4543));
   CLKBUFX2TS FE_OFC276_n4543 (.Y(FE_OFN276_n4543), 
	.A(FE_OFN273_n4543));
   CLKBUFX2TS FE_OFC275_n4543 (.Y(FE_OFN275_n4543), 
	.A(FE_OFN271_n4543));
   CLKBUFX2TS FE_OFC274_n4543 (.Y(FE_OFN274_n4543), 
	.A(FE_OFN273_n4543));
   CLKBUFX2TS FE_OFC273_n4543 (.Y(FE_OFN273_n4543), 
	.A(FE_OFN270_n4543));
   CLKBUFX2TS FE_OFC272_n4543 (.Y(FE_OFN272_n4543), 
	.A(FE_OFN268_n4543));
   CLKBUFX2TS FE_OFC271_n4543 (.Y(FE_OFN271_n4543), 
	.A(FE_OFN269_n4543));
   CLKBUFX2TS FE_OFC270_n4543 (.Y(FE_OFN270_n4543), 
	.A(FE_OFN269_n4543));
   CLKBUFX2TS FE_OFC269_n4543 (.Y(FE_OFN269_n4543), 
	.A(FE_OFN267_n4543));
   CLKBUFX2TS FE_OFC268_n4543 (.Y(FE_OFN268_n4543), 
	.A(FE_OFN266_n4543));
   CLKBUFX2TS FE_OFC267_n4543 (.Y(FE_OFN267_n4543), 
	.A(FE_OFN266_n4543));
   CLKBUFX2TS FE_OFC266_n4543 (.Y(FE_OFN266_n4543), 
	.A(n4543));
   CLKBUFX2TS FE_OFC265_n4544 (.Y(FE_OFN265_n4544), 
	.A(FE_OFN264_n4544));
   CLKBUFX2TS FE_OFC264_n4544 (.Y(FE_OFN264_n4544), 
	.A(FE_OFN263_n4544));
   CLKBUFX2TS FE_OFC263_n4544 (.Y(FE_OFN263_n4544), 
	.A(FE_OFN262_n4544));
   CLKBUFX2TS FE_OFC262_n4544 (.Y(FE_OFN262_n4544), 
	.A(FE_OFN259_n4544));
   CLKBUFX2TS FE_OFC261_n4544 (.Y(FE_OFN261_n4544), 
	.A(FE_OFN260_n4544));
   CLKBUFX2TS FE_OFC260_n4544 (.Y(FE_OFN260_n4544), 
	.A(FE_OFN257_n4544));
   CLKBUFX2TS FE_OFC259_n4544 (.Y(FE_OFN259_n4544), 
	.A(FE_OFN258_n4544));
   CLKBUFX2TS FE_OFC258_n4544 (.Y(FE_OFN258_n4544), 
	.A(FE_OFN256_n4544));
   CLKBUFX2TS FE_OFC257_n4544 (.Y(FE_OFN257_n4544), 
	.A(n4544));
   CLKBUFX2TS FE_OFC256_n4544 (.Y(FE_OFN256_n4544), 
	.A(n4544));
   CLKBUFX2TS FE_OFC255_n4537 (.Y(FE_OFN255_n4537), 
	.A(FE_OFN254_n4537));
   CLKBUFX2TS FE_OFC254_n4537 (.Y(FE_OFN254_n4537), 
	.A(FE_OFN253_n4537));
   CLKBUFX2TS FE_OFC253_n4537 (.Y(FE_OFN253_n4537), 
	.A(FE_OFN252_n4537));
   CLKBUFX2TS FE_OFC252_n4537 (.Y(FE_OFN252_n4537), 
	.A(FE_OFN251_n4537));
   CLKBUFX2TS FE_OFC251_n4537 (.Y(FE_OFN251_n4537), 
	.A(FE_OFN248_n4537));
   CLKBUFX2TS FE_OFC250_n4537 (.Y(FE_OFN250_n4537), 
	.A(FE_OFN248_n4537));
   CLKBUFX2TS FE_OFC249_n4537 (.Y(FE_OFN249_n4537), 
	.A(FE_OFN246_n4537));
   CLKBUFX2TS FE_OFC248_n4537 (.Y(FE_OFN248_n4537), 
	.A(FE_OFN245_n4537));
   CLKBUFX2TS FE_OFC247_n4537 (.Y(FE_OFN247_n4537), 
	.A(FE_OFN245_n4537));
   CLKBUFX2TS FE_OFC246_n4537 (.Y(FE_OFN246_n4537), 
	.A(FE_OFN244_n4537));
   CLKBUFX2TS FE_OFC245_n4537 (.Y(FE_OFN245_n4537), 
	.A(n4537));
   CLKBUFX2TS FE_OFC244_n4537 (.Y(FE_OFN244_n4537), 
	.A(n4537));
   CLKBUFX2TS FE_OFC243_n4531 (.Y(FE_OFN243_n4531), 
	.A(FE_OFN242_n4531));
   CLKBUFX2TS FE_OFC242_n4531 (.Y(FE_OFN242_n4531), 
	.A(FE_OFN238_n4531));
   CLKBUFX2TS FE_OFC241_n4531 (.Y(FE_OFN241_n4531), 
	.A(FE_OFN239_n4531));
   CLKBUFX2TS FE_OFC240_n4531 (.Y(FE_OFN240_n4531), 
	.A(FE_OFN239_n4531));
   CLKBUFX2TS FE_OFC239_n4531 (.Y(FE_OFN239_n4531), 
	.A(FE_OFN236_n4531));
   CLKBUFX2TS FE_OFC238_n4531 (.Y(FE_OFN238_n4531), 
	.A(FE_OFN236_n4531));
   CLKBUFX2TS FE_OFC237_n4531 (.Y(FE_OFN237_n4531), 
	.A(FE_OFN234_n4531));
   CLKBUFX2TS FE_OFC236_n4531 (.Y(FE_OFN236_n4531), 
	.A(FE_OFN235_n4531));
   CLKBUFX2TS FE_OFC235_n4531 (.Y(FE_OFN235_n4531), 
	.A(FE_OFN233_n4531));
   CLKBUFX2TS FE_OFC234_n4531 (.Y(FE_OFN234_n4531), 
	.A(FE_OFN232_n4531));
   CLKBUFX2TS FE_OFC233_n4531 (.Y(FE_OFN233_n4531), 
	.A(n4531));
   CLKBUFX2TS FE_OFC232_n4531 (.Y(FE_OFN232_n4531), 
	.A(n4531));
   CLKBUFX2TS FE_OFC231_n4525 (.Y(FE_OFN231_n4525), 
	.A(FE_OFN230_n4525));
   CLKBUFX2TS FE_OFC230_n4525 (.Y(FE_OFN230_n4525), 
	.A(FE_OFN229_n4525));
   CLKBUFX2TS FE_OFC229_n4525 (.Y(FE_OFN229_n4525), 
	.A(FE_OFN227_n4525));
   CLKBUFX2TS FE_OFC228_n4525 (.Y(FE_OFN228_n4525), 
	.A(FE_OFN227_n4525));
   CLKBUFX2TS FE_OFC227_n4525 (.Y(FE_OFN227_n4525), 
	.A(FE_OFN225_n4525));
   CLKBUFX2TS FE_OFC226_n4525 (.Y(FE_OFN226_n4525), 
	.A(FE_OFN223_n4525));
   CLKBUFX2TS FE_OFC225_n4525 (.Y(FE_OFN225_n4525), 
	.A(FE_OFN223_n4525));
   CLKBUFX2TS FE_OFC224_n4525 (.Y(FE_OFN224_n4525), 
	.A(FE_OFN222_n4525));
   CLKBUFX2TS FE_OFC223_n4525 (.Y(FE_OFN223_n4525), 
	.A(FE_OFN222_n4525));
   CLKBUFX2TS FE_OFC222_n4525 (.Y(FE_OFN222_n4525), 
	.A(FE_OFN221_n4525));
   CLKBUFX2TS FE_OFC221_n4525 (.Y(FE_OFN221_n4525), 
	.A(n4525));
   CLKBUFX2TS FE_OFC220_n4519 (.Y(FE_OFN220_n4519), 
	.A(FE_OFN219_n4519));
   CLKBUFX2TS FE_OFC219_n4519 (.Y(FE_OFN219_n4519), 
	.A(FE_OFN216_n4519));
   CLKBUFX2TS FE_OFC218_n4519 (.Y(FE_OFN218_n4519), 
	.A(FE_OFN215_n4519));
   CLKBUFX2TS FE_OFC217_n4519 (.Y(FE_OFN217_n4519), 
	.A(FE_OFN215_n4519));
   CLKBUFX2TS FE_OFC216_n4519 (.Y(FE_OFN216_n4519), 
	.A(FE_OFN214_n4519));
   CLKBUFX2TS FE_OFC215_n4519 (.Y(FE_OFN215_n4519), 
	.A(FE_OFN213_n4519));
   CLKBUFX2TS FE_OFC214_n4519 (.Y(FE_OFN214_n4519), 
	.A(FE_OFN211_n4519));
   CLKBUFX2TS FE_OFC213_n4519 (.Y(FE_OFN213_n4519), 
	.A(FE_OFN212_n4519));
   CLKBUFX2TS FE_OFC212_n4519 (.Y(FE_OFN212_n4519), 
	.A(FE_OFN210_n4519));
   CLKBUFX2TS FE_OFC211_n4519 (.Y(FE_OFN211_n4519), 
	.A(FE_OFN210_n4519));
   CLKBUFX2TS FE_OFC210_n4519 (.Y(FE_OFN210_n4519), 
	.A(n4519));
   CLKBUFX2TS FE_OFC209_n4519 (.Y(FE_OFN209_n4519), 
	.A(n4519));
   CLKBUFX2TS FE_OFC208_n4513 (.Y(FE_OFN208_n4513), 
	.A(FE_OFN207_n4513));
   CLKBUFX2TS FE_OFC207_n4513 (.Y(FE_OFN207_n4513), 
	.A(FE_OFN204_n4513));
   CLKBUFX2TS FE_OFC206_n4513 (.Y(FE_OFN206_n4513), 
	.A(FE_OFN203_n4513));
   CLKBUFX2TS FE_OFC205_n4513 (.Y(FE_OFN205_n4513), 
	.A(FE_OFN203_n4513));
   CLKBUFX2TS FE_OFC204_n4513 (.Y(FE_OFN204_n4513), 
	.A(FE_OFN201_n4513));
   CLKBUFX2TS FE_OFC203_n4513 (.Y(FE_OFN203_n4513), 
	.A(FE_OFN202_n4513));
   CLKBUFX2TS FE_OFC202_n4513 (.Y(FE_OFN202_n4513), 
	.A(FE_OFN200_n4513));
   CLKBUFX2TS FE_OFC201_n4513 (.Y(FE_OFN201_n4513), 
	.A(FE_OFN200_n4513));
   CLKBUFX2TS FE_OFC200_n4513 (.Y(FE_OFN200_n4513), 
	.A(FE_OFN197_n4513));
   CLKBUFX2TS FE_OFC199_n4513 (.Y(FE_OFN199_n4513), 
	.A(FE_OFN198_n4513));
   CLKBUFX2TS FE_OFC198_n4513 (.Y(FE_OFN198_n4513), 
	.A(n4513));
   CLKBUFX2TS FE_OFC197_n4513 (.Y(FE_OFN197_n4513), 
	.A(n4513));
   CLKBUFX2TS FE_OFC196_n4514 (.Y(FE_OFN196_n4514), 
	.A(FE_OFN195_n4514));
   CLKBUFX2TS FE_OFC195_n4514 (.Y(FE_OFN195_n4514), 
	.A(FE_OFN192_n4514));
   CLKBUFX2TS FE_OFC194_n4514 (.Y(FE_OFN194_n4514), 
	.A(FE_OFN193_n4514));
   CLKBUFX2TS FE_OFC193_n4514 (.Y(FE_OFN193_n4514), 
	.A(FE_OFN190_n4514));
   CLKBUFX2TS FE_OFC192_n4514 (.Y(FE_OFN192_n4514), 
	.A(FE_OFN191_n4514));
   CLKBUFX2TS FE_OFC191_n4514 (.Y(FE_OFN191_n4514), 
	.A(FE_OFN189_n4514));
   CLKBUFX2TS FE_OFC190_n4514 (.Y(FE_OFN190_n4514), 
	.A(FE_OFN188_n4514));
   CLKBUFX2TS FE_OFC189_n4514 (.Y(FE_OFN189_n4514), 
	.A(FE_OFN187_n4514));
   CLKBUFX2TS FE_OFC188_n4514 (.Y(FE_OFN188_n4514), 
	.A(n4514));
   CLKBUFX2TS FE_OFC187_n4514 (.Y(FE_OFN187_n4514), 
	.A(n4514));
   CLKBUFX2TS FE_OFC186_n4507 (.Y(FE_OFN186_n4507), 
	.A(FE_OFN185_n4507));
   CLKBUFX2TS FE_OFC185_n4507 (.Y(FE_OFN185_n4507), 
	.A(FE_OFN184_n4507));
   CLKBUFX2TS FE_OFC184_n4507 (.Y(FE_OFN184_n4507), 
	.A(FE_OFN182_n4507));
   CLKBUFX2TS FE_OFC183_n4507 (.Y(FE_OFN183_n4507), 
	.A(FE_OFN181_n4507));
   CLKBUFX2TS FE_OFC182_n4507 (.Y(FE_OFN182_n4507), 
	.A(FE_OFN179_n4507));
   CLKBUFX2TS FE_OFC181_n4507 (.Y(FE_OFN181_n4507), 
	.A(FE_OFN180_n4507));
   CLKBUFX2TS FE_OFC180_n4507 (.Y(FE_OFN180_n4507), 
	.A(FE_OFN177_n4507));
   CLKBUFX2TS FE_OFC179_n4507 (.Y(FE_OFN179_n4507), 
	.A(FE_OFN178_n4507));
   CLKBUFX2TS FE_OFC178_n4507 (.Y(FE_OFN178_n4507), 
	.A(FE_OFN176_n4507));
   CLKBUFX2TS FE_OFC177_n4507 (.Y(FE_OFN177_n4507), 
	.A(FE_OFN176_n4507));
   CLKBUFX2TS FE_OFC176_n4507 (.Y(FE_OFN176_n4507), 
	.A(FE_OFN175_n4507));
   CLKBUFX2TS FE_OFC175_n4507 (.Y(FE_OFN175_n4507), 
	.A(n4507));
   CLKBUFX2TS FE_OFC174_n8054 (.Y(FE_OFN174_n8054), 
	.A(FE_OFN173_n8054));
   CLKBUFX2TS FE_OFC173_n8054 (.Y(FE_OFN173_n8054), 
	.A(n8054));
   CLKBUFX2TS FE_OFC172_n4495 (.Y(FE_OFN172_n4495), 
	.A(FE_OFN171_n4495));
   CLKBUFX2TS FE_OFC171_n4495 (.Y(FE_OFN171_n4495), 
	.A(FE_OFN170_n4495));
   CLKBUFX2TS FE_OFC170_n4495 (.Y(FE_OFN170_n4495), 
	.A(FE_OFN168_n4495));
   CLKBUFX2TS FE_OFC169_n4495 (.Y(FE_OFN169_n4495), 
	.A(FE_OFN167_n4495));
   CLKBUFX2TS FE_OFC168_n4495 (.Y(FE_OFN168_n4495), 
	.A(FE_OFN166_n4495));
   CLKBUFX2TS FE_OFC167_n4495 (.Y(FE_OFN167_n4495), 
	.A(FE_OFN165_n4495));
   CLKBUFX2TS FE_OFC166_n4495 (.Y(FE_OFN166_n4495), 
	.A(FE_OFN164_n4495));
   CLKBUFX2TS FE_OFC165_n4495 (.Y(FE_OFN165_n4495), 
	.A(FE_OFN163_n4495));
   CLKBUFX2TS FE_OFC164_n4495 (.Y(FE_OFN164_n4495), 
	.A(FE_OFN163_n4495));
   CLKBUFX2TS FE_OFC163_n4495 (.Y(FE_OFN163_n4495), 
	.A(FE_OFN162_n4495));
   CLKBUFX2TS FE_OFC162_n4495 (.Y(FE_OFN162_n4495), 
	.A(FE_OFN161_n4495));
   CLKBUFX2TS FE_OFC161_n4495 (.Y(FE_OFN161_n4495), 
	.A(n4495));
   CLKBUFX2TS FE_OFC160_n4496 (.Y(FE_OFN160_n4496), 
	.A(FE_OFN157_n4496));
   CLKBUFX2TS FE_OFC159_n4496 (.Y(FE_OFN159_n4496), 
	.A(FE_OFN156_n4496));
   CLKBUFX2TS FE_OFC158_n4496 (.Y(FE_OFN158_n4496), 
	.A(FE_OFN156_n4496));
   CLKBUFX2TS FE_OFC157_n4496 (.Y(FE_OFN157_n4496), 
	.A(FE_OFN155_n4496));
   CLKBUFX2TS FE_OFC156_n4496 (.Y(FE_OFN156_n4496), 
	.A(FE_OFN154_n4496));
   CLKBUFX2TS FE_OFC155_n4496 (.Y(FE_OFN155_n4496), 
	.A(FE_OFN153_n4496));
   CLKBUFX2TS FE_OFC154_n4496 (.Y(FE_OFN154_n4496), 
	.A(FE_OFN152_n4496));
   CLKBUFX2TS FE_OFC153_n4496 (.Y(FE_OFN153_n4496), 
	.A(FE_OFN152_n4496));
   CLKBUFX2TS FE_OFC152_n4496 (.Y(FE_OFN152_n4496), 
	.A(FE_OFN151_n4496));
   CLKBUFX2TS FE_OFC151_n4496 (.Y(FE_OFN151_n4496), 
	.A(n4496));
   CLKBUFX2TS FE_OFC150_n4489 (.Y(FE_OFN150_n4489), 
	.A(FE_OFN149_n4489));
   CLKBUFX2TS FE_OFC149_n4489 (.Y(FE_OFN149_n4489), 
	.A(FE_OFN148_n4489));
   CLKBUFX2TS FE_OFC148_n4489 (.Y(FE_OFN148_n4489), 
	.A(FE_OFN147_n4489));
   CLKBUFX2TS FE_OFC147_n4489 (.Y(FE_OFN147_n4489), 
	.A(FE_OFN146_n4489));
   CLKBUFX2TS FE_OFC146_n4489 (.Y(FE_OFN146_n4489), 
	.A(FE_OFN144_n4489));
   CLKBUFX2TS FE_OFC145_n4489 (.Y(FE_OFN145_n4489), 
	.A(FE_OFN143_n4489));
   CLKBUFX2TS FE_OFC144_n4489 (.Y(FE_OFN144_n4489), 
	.A(FE_OFN141_n4489));
   CLKBUFX2TS FE_OFC143_n4489 (.Y(FE_OFN143_n4489), 
	.A(FE_OFN142_n4489));
   CLKBUFX2TS FE_OFC142_n4489 (.Y(FE_OFN142_n4489), 
	.A(FE_OFN140_n4489));
   CLKBUFX2TS FE_OFC141_n4489 (.Y(FE_OFN141_n4489), 
	.A(FE_OFN140_n4489));
   CLKBUFX2TS FE_OFC140_n4489 (.Y(FE_OFN140_n4489), 
	.A(FE_OFN139_n4489));
   CLKBUFX2TS FE_OFC139_n4489 (.Y(FE_OFN139_n4489), 
	.A(n4489));
   CLKBUFX2TS FE_OFC138_n4490 (.Y(FE_OFN138_n4490), 
	.A(FE_OFN137_n4490));
   CLKBUFX2TS FE_OFC137_n4490 (.Y(FE_OFN137_n4490), 
	.A(FE_OFN136_n4490));
   CLKBUFX2TS FE_OFC136_n4490 (.Y(FE_OFN136_n4490), 
	.A(FE_OFN135_n4490));
   CLKBUFX2TS FE_OFC135_n4490 (.Y(FE_OFN135_n4490), 
	.A(FE_OFN134_n4490));
   CLKBUFX2TS FE_OFC134_n4490 (.Y(FE_OFN134_n4490), 
	.A(FE_OFN132_n4490));
   CLKBUFX2TS FE_OFC133_n4490 (.Y(FE_OFN133_n4490), 
	.A(FE_OFN131_n4490));
   CLKBUFX2TS FE_OFC132_n4490 (.Y(FE_OFN132_n4490), 
	.A(FE_OFN131_n4490));
   CLKBUFX2TS FE_OFC131_n4490 (.Y(FE_OFN131_n4490), 
	.A(FE_OFN130_n4490));
   CLKBUFX2TS FE_OFC130_n4490 (.Y(FE_OFN130_n4490), 
	.A(FE_OFN129_n4490));
   CLKBUFX2TS FE_OFC129_n4490 (.Y(FE_OFN129_n4490), 
	.A(n4490));
   CLKBUFX2TS FE_OFC128_n4502 (.Y(FE_OFN128_n4502), 
	.A(FE_OFN127_n4502));
   CLKBUFX2TS FE_OFC127_n4502 (.Y(FE_OFN127_n4502), 
	.A(FE_OFN126_n4502));
   CLKBUFX2TS FE_OFC126_n4502 (.Y(FE_OFN126_n4502), 
	.A(FE_OFN125_n4502));
   CLKBUFX2TS FE_OFC125_n4502 (.Y(FE_OFN125_n4502), 
	.A(FE_OFN123_n4502));
   CLKINVX1TS FE_OFC124_n4502 (.Y(FE_OFN124_n4502), 
	.A(FE_OFN121_n4502));
   CLKINVX1TS FE_OFC123_n4502 (.Y(FE_OFN123_n4502), 
	.A(FE_OFN121_n4502));
   CLKBUFX2TS FE_OFC122_n4502 (.Y(FE_OFN122_n4502), 
	.A(FE_OFN119_n4502));
   CLKINVX1TS FE_OFC121_n4502 (.Y(FE_OFN121_n4502), 
	.A(FE_OFN116_n4502));
   CLKINVX1TS FE_OFC120_n4502 (.Y(FE_OFN120_n4502), 
	.A(FE_OFN117_n4502));
   CLKINVX1TS FE_OFC119_n4502 (.Y(FE_OFN119_n4502), 
	.A(FE_OFN117_n4502));
   CLKBUFX2TS FE_OFC118_n4502 (.Y(FE_OFN118_n4502), 
	.A(FE_OFN116_n4502));
   CLKINVX1TS FE_OFC117_n4502 (.Y(FE_OFN117_n4502), 
	.A(FE_OFN115_n4502));
   CLKBUFX2TS FE_OFC116_n4502 (.Y(FE_OFN116_n4502), 
	.A(FE_OFN115_n4502));
   CLKBUFX2TS FE_OFC115_n4502 (.Y(FE_OFN115_n4502), 
	.A(n4502));
   CLKBUFX2TS FE_OFC114_n4508 (.Y(FE_OFN114_n4508), 
	.A(FE_OFN113_n4508));
   CLKBUFX2TS FE_OFC113_n4508 (.Y(FE_OFN113_n4508), 
	.A(FE_OFN111_n4508));
   CLKBUFX2TS FE_OFC112_n4508 (.Y(FE_OFN112_n4508), 
	.A(FE_OFN110_n4508));
   CLKBUFX2TS FE_OFC111_n4508 (.Y(FE_OFN111_n4508), 
	.A(FE_OFN109_n4508));
   CLKBUFX2TS FE_OFC110_n4508 (.Y(FE_OFN110_n4508), 
	.A(FE_OFN108_n4508));
   CLKBUFX2TS FE_OFC109_n4508 (.Y(FE_OFN109_n4508), 
	.A(FE_OFN107_n4508));
   CLKBUFX2TS FE_OFC108_n4508 (.Y(FE_OFN108_n4508), 
	.A(FE_OFN106_n4508));
   CLKBUFX2TS FE_OFC107_n4508 (.Y(FE_OFN107_n4508), 
	.A(FE_OFN105_n4508));
   CLKBUFX2TS FE_OFC106_n4508 (.Y(FE_OFN106_n4508), 
	.A(n4508));
   CLKBUFX2TS FE_OFC105_n4508 (.Y(FE_OFN105_n4508), 
	.A(n4508));
   CLKBUFX2TS FE_OFC104_n4520 (.Y(FE_OFN104_n4520), 
	.A(FE_OFN103_n4520));
   CLKBUFX2TS FE_OFC103_n4520 (.Y(FE_OFN103_n4520), 
	.A(FE_OFN102_n4520));
   CLKBUFX2TS FE_OFC102_n4520 (.Y(FE_OFN102_n4520), 
	.A(FE_OFN99_n4520));
   CLKBUFX2TS FE_OFC101_n4520 (.Y(FE_OFN101_n4520), 
	.A(FE_OFN98_n4520));
   CLKBUFX2TS FE_OFC100_n4520 (.Y(FE_OFN100_n4520), 
	.A(FE_OFN98_n4520));
   CLKBUFX2TS FE_OFC99_n4520 (.Y(FE_OFN99_n4520), 
	.A(FE_OFN96_n4520));
   CLKBUFX2TS FE_OFC98_n4520 (.Y(FE_OFN98_n4520), 
	.A(FE_OFN95_n4520));
   CLKBUFX2TS FE_OFC97_n4520 (.Y(FE_OFN97_n4520), 
	.A(FE_OFN95_n4520));
   CLKBUFX2TS FE_OFC96_n4520 (.Y(FE_OFN96_n4520), 
	.A(n4520));
   CLKBUFX2TS FE_OFC95_n4520 (.Y(FE_OFN95_n4520), 
	.A(n4520));
   CLKBUFX2TS FE_OFC94_n4526 (.Y(FE_OFN94_n4526), 
	.A(FE_OFN93_n4526));
   CLKBUFX2TS FE_OFC93_n4526 (.Y(FE_OFN93_n4526), 
	.A(FE_OFN92_n4526));
   CLKBUFX2TS FE_OFC92_n4526 (.Y(FE_OFN92_n4526), 
	.A(FE_OFN91_n4526));
   CLKBUFX2TS FE_OFC91_n4526 (.Y(FE_OFN91_n4526), 
	.A(FE_OFN90_n4526));
   CLKBUFX2TS FE_OFC90_n4526 (.Y(FE_OFN90_n4526), 
	.A(FE_OFN87_n4526));
   CLKBUFX2TS FE_OFC89_n4526 (.Y(FE_OFN89_n4526), 
	.A(FE_OFN86_n4526));
   CLKBUFX2TS FE_OFC88_n4526 (.Y(FE_OFN88_n4526), 
	.A(FE_OFN86_n4526));
   CLKBUFX2TS FE_OFC87_n4526 (.Y(FE_OFN87_n4526), 
	.A(FE_OFN84_n4526));
   CLKBUFX2TS FE_OFC86_n4526 (.Y(FE_OFN86_n4526), 
	.A(FE_OFN84_n4526));
   CLKBUFX2TS FE_OFC85_n4526 (.Y(FE_OFN85_n4526), 
	.A(n4526));
   CLKBUFX2TS FE_OFC84_n4526 (.Y(FE_OFN84_n4526), 
	.A(n4526));
   CLKBUFX2TS FE_OFC83_n3796 (.Y(FE_OFN83_n3796), 
	.A(FE_OFN81_n3796));
   CLKBUFX2TS FE_OFC82_n3796 (.Y(FE_OFN82_n3796), 
	.A(FE_OFN80_n3796));
   CLKBUFX2TS FE_OFC81_n3796 (.Y(FE_OFN81_n3796), 
	.A(FE_OFN79_n3796));
   CLKBUFX2TS FE_OFC80_n3796 (.Y(FE_OFN80_n3796), 
	.A(FE_OFN78_n3796));
   CLKBUFX2TS FE_OFC79_n3796 (.Y(FE_OFN79_n3796), 
	.A(FE_OFN77_n3796));
   CLKBUFX2TS FE_OFC78_n3796 (.Y(FE_OFN78_n3796), 
	.A(FE_OFN76_n3796));
   CLKBUFX2TS FE_OFC77_n3796 (.Y(FE_OFN77_n3796), 
	.A(FE_OFN75_n3796));
   CLKBUFX2TS FE_OFC76_n3796 (.Y(FE_OFN76_n3796), 
	.A(FE_OFN75_n3796));
   CLKBUFX2TS FE_OFC75_n3796 (.Y(FE_OFN75_n3796), 
	.A(FE_OFN74_n3796));
   CLKBUFX2TS FE_OFC74_n3796 (.Y(FE_OFN74_n3796), 
	.A(FE_OFN73_n3796));
   CLKBUFX2TS FE_OFC73_n3796 (.Y(FE_OFN73_n3796), 
	.A(n3796));
   CLKBUFX2TS FE_OFC72_n3797 (.Y(FE_OFN72_n3797), 
	.A(FE_OFN70_n3797));
   CLKBUFX2TS FE_OFC71_n3797 (.Y(FE_OFN71_n3797), 
	.A(FE_OFN69_n3797));
   CLKBUFX2TS FE_OFC70_n3797 (.Y(FE_OFN70_n3797), 
	.A(FE_OFN68_n3797));
   CLKBUFX2TS FE_OFC69_n3797 (.Y(FE_OFN69_n3797), 
	.A(FE_OFN67_n3797));
   CLKBUFX2TS FE_OFC68_n3797 (.Y(FE_OFN68_n3797), 
	.A(FE_OFN66_n3797));
   CLKBUFX2TS FE_OFC67_n3797 (.Y(FE_OFN67_n3797), 
	.A(FE_OFN65_n3797));
   CLKBUFX2TS FE_OFC66_n3797 (.Y(FE_OFN66_n3797), 
	.A(FE_OFN64_n3797));
   CLKBUFX2TS FE_OFC65_n3797 (.Y(FE_OFN65_n3797), 
	.A(FE_OFN64_n3797));
   CLKBUFX2TS FE_OFC64_n3797 (.Y(FE_OFN64_n3797), 
	.A(FE_OFN63_n3797));
   CLKBUFX2TS FE_OFC63_n3797 (.Y(FE_OFN63_n3797), 
	.A(n3797));
   CLKBUFX2TS FE_OFC62_n4532 (.Y(FE_OFN62_n4532), 
	.A(FE_OFN61_n4532));
   CLKBUFX2TS FE_OFC61_n4532 (.Y(FE_OFN61_n4532), 
	.A(FE_OFN58_n4532));
   CLKBUFX2TS FE_OFC60_n4532 (.Y(FE_OFN60_n4532), 
	.A(FE_OFN57_n4532));
   CLKBUFX2TS FE_OFC59_n4532 (.Y(FE_OFN59_n4532), 
	.A(FE_OFN56_n4532));
   CLKBUFX2TS FE_OFC58_n4532 (.Y(FE_OFN58_n4532), 
	.A(FE_OFN55_n4532));
   CLKBUFX2TS FE_OFC57_n4532 (.Y(FE_OFN57_n4532), 
	.A(FE_OFN55_n4532));
   CLKBUFX2TS FE_OFC56_n4532 (.Y(FE_OFN56_n4532), 
	.A(FE_OFN54_n4532));
   CLKBUFX2TS FE_OFC55_n4532 (.Y(FE_OFN55_n4532), 
	.A(FE_OFN53_n4532));
   CLKBUFX2TS FE_OFC54_n4532 (.Y(FE_OFN54_n4532), 
	.A(FE_OFN53_n4532));
   CLKBUFX2TS FE_OFC53_n4532 (.Y(FE_OFN53_n4532), 
	.A(n4532));
   CLKBUFX2TS FE_OFC52_n4538 (.Y(FE_OFN52_n4538), 
	.A(FE_OFN51_n4538));
   CLKBUFX2TS FE_OFC51_n4538 (.Y(FE_OFN51_n4538), 
	.A(FE_OFN49_n4538));
   CLKBUFX2TS FE_OFC50_n4538 (.Y(FE_OFN50_n4538), 
	.A(FE_OFN48_n4538));
   CLKBUFX2TS FE_OFC49_n4538 (.Y(FE_OFN49_n4538), 
	.A(FE_OFN47_n4538));
   CLKBUFX2TS FE_OFC48_n4538 (.Y(FE_OFN48_n4538), 
	.A(FE_OFN46_n4538));
   CLKBUFX2TS FE_OFC47_n4538 (.Y(FE_OFN47_n4538), 
	.A(FE_OFN45_n4538));
   CLKBUFX2TS FE_OFC46_n4538 (.Y(FE_OFN46_n4538), 
	.A(FE_OFN43_n4538));
   CLKBUFX2TS FE_OFC45_n4538 (.Y(FE_OFN45_n4538), 
	.A(FE_OFN44_n4538));
   CLKBUFX2TS FE_OFC44_n4538 (.Y(FE_OFN44_n4538), 
	.A(n4538));
   CLKBUFX2TS FE_OFC43_n4538 (.Y(FE_OFN43_n4538), 
	.A(n4538));
   CLKBUFX2TS FE_OFC42_n4550 (.Y(FE_OFN42_n4550), 
	.A(FE_OFN40_n4550));
   CLKBUFX2TS FE_OFC41_n4550 (.Y(FE_OFN41_n4550), 
	.A(FE_OFN40_n4550));
   CLKBUFX2TS FE_OFC40_n4550 (.Y(FE_OFN40_n4550), 
	.A(FE_OFN39_n4550));
   CLKBUFX2TS FE_OFC39_n4550 (.Y(FE_OFN39_n4550), 
	.A(FE_OFN38_n4550));
   CLKBUFX2TS FE_OFC38_n4550 (.Y(FE_OFN38_n4550), 
	.A(FE_OFN37_n4550));
   CLKBUFX2TS FE_OFC37_n4550 (.Y(FE_OFN37_n4550), 
	.A(FE_OFN36_n4550));
   CLKBUFX2TS FE_OFC36_n4550 (.Y(FE_OFN36_n4550), 
	.A(FE_OFN35_n4550));
   CLKBUFX2TS FE_OFC35_n4550 (.Y(FE_OFN35_n4550), 
	.A(FE_OFN34_n4550));
   CLKBUFX2TS FE_OFC34_n4550 (.Y(FE_OFN34_n4550), 
	.A(FE_OFN33_n4550));
   CLKBUFX2TS FE_OFC33_n4550 (.Y(FE_OFN33_n4550), 
	.A(n4550));
   CLKBUFX2TS FE_OFC32_n4562 (.Y(FE_OFN32_n4562), 
	.A(FE_OFN30_n4562));
   CLKBUFX2TS FE_OFC31_n4562 (.Y(FE_OFN31_n4562), 
	.A(FE_OFN30_n4562));
   CLKBUFX2TS FE_OFC30_n4562 (.Y(FE_OFN30_n4562), 
	.A(FE_OFN29_n4562));
   CLKBUFX2TS FE_OFC29_n4562 (.Y(FE_OFN29_n4562), 
	.A(FE_OFN27_n4562));
   CLKBUFX2TS FE_OFC28_n4562 (.Y(FE_OFN28_n4562), 
	.A(FE_OFN26_n4562));
   CLKBUFX2TS FE_OFC27_n4562 (.Y(FE_OFN27_n4562), 
	.A(FE_OFN26_n4562));
   CLKBUFX2TS FE_OFC26_n4562 (.Y(FE_OFN26_n4562), 
	.A(FE_OFN23_n4562));
   CLKBUFX2TS FE_OFC25_n4562 (.Y(FE_OFN25_n4562), 
	.A(FE_OFN24_n4562));
   CLKBUFX2TS FE_OFC24_n4562 (.Y(FE_OFN24_n4562), 
	.A(FE_OFN22_n4562));
   CLKBUFX2TS FE_OFC23_n4562 (.Y(FE_OFN23_n4562), 
	.A(n4562));
   CLKBUFX2TS FE_OFC22_n4562 (.Y(FE_OFN22_n4562), 
	.A(n4562));
   CLKBUFX2TS FE_OFC21_n4568 (.Y(FE_OFN21_n4568), 
	.A(FE_OFN20_n4568));
   CLKBUFX2TS FE_OFC20_n4568 (.Y(FE_OFN20_n4568), 
	.A(FE_OFN18_n4568));
   CLKBUFX2TS FE_OFC19_n4568 (.Y(FE_OFN19_n4568), 
	.A(FE_OFN17_n4568));
   CLKBUFX2TS FE_OFC18_n4568 (.Y(FE_OFN18_n4568), 
	.A(FE_OFN17_n4568));
   CLKBUFX2TS FE_OFC17_n4568 (.Y(FE_OFN17_n4568), 
	.A(FE_OFN16_n4568));
   CLKBUFX2TS FE_OFC16_n4568 (.Y(FE_OFN16_n4568), 
	.A(FE_OFN15_n4568));
   CLKBUFX2TS FE_OFC15_n4568 (.Y(FE_OFN15_n4568), 
	.A(FE_OFN13_n4568));
   CLKINVX1TS FE_OFC14_n4568 (.Y(FE_OFN14_n4568), 
	.A(FE_OFN12_n4568));
   CLKINVX1TS FE_OFC13_n4568 (.Y(FE_OFN13_n4568), 
	.A(FE_OFN12_n4568));
   CLKINVX1TS FE_OFC12_n4568 (.Y(FE_OFN12_n4568), 
	.A(FE_OFN11_n4568));
   CLKBUFX2TS FE_OFC11_n4568 (.Y(FE_OFN11_n4568), 
	.A(FE_OFN10_n4568));
   CLKBUFX2TS FE_OFC10_n4568 (.Y(FE_OFN10_n4568), 
	.A(n4568));
   CLKBUFX2TS FE_OFC9_n4574 (.Y(FE_OFN9_n4574), 
	.A(FE_OFN8_n4574));
   CLKBUFX2TS FE_OFC8_n4574 (.Y(FE_OFN8_n4574), 
	.A(FE_OFN7_n4574));
   CLKBUFX2TS FE_OFC7_n4574 (.Y(FE_OFN7_n4574), 
	.A(FE_OFN6_n4574));
   CLKBUFX2TS FE_OFC6_n4574 (.Y(FE_OFN6_n4574), 
	.A(FE_OFN5_n4574));
   CLKBUFX2TS FE_OFC5_n4574 (.Y(FE_OFN5_n4574), 
	.A(FE_OFN4_n4574));
   CLKBUFX2TS FE_OFC4_n4574 (.Y(FE_OFN4_n4574), 
	.A(FE_OFN3_n4574));
   CLKBUFX2TS FE_OFC3_n4574 (.Y(FE_OFN3_n4574), 
	.A(FE_OFN2_n4574));
   CLKBUFX2TS FE_OFC2_n4574 (.Y(FE_OFN2_n4574), 
	.A(FE_OFN1_n4574));
   CLKBUFX2TS FE_OFC1_n4574 (.Y(FE_OFN1_n4574), 
	.A(FE_OFN0_n4574));
   CLKBUFX2TS FE_OFC0_n4574 (.Y(FE_OFN0_n4574), 
	.A(n4574));
   BUFX2TS FE_MDBC14_U5721 (.Y(FE_MDBN14_), 
	.A(fft_data_in[31]));
   BUFX2TS FE_MDBC13_U5679 (.Y(FE_MDBN13_), 
	.A(fft_data_in[30]));
   BUFX2TS FE_MDBC12_U5586 (.Y(FE_MDBN12_), 
	.A(fft_data_in[29]));
   BUFX2TS FE_MDBC11_U5490 (.Y(FE_MDBN11_), 
	.A(fft_data_in[28]));
   BUFX2TS FE_MDBC10_U5445 (.Y(FE_MDBN10_), 
	.A(fft_data_in[27]));
   BUFX2TS FE_MDBC9_U5223 (.Y(FE_MDBN9_), 
	.A(fft_data_in[26]));
   BUFX2TS FE_MDBC8_U5221 (.Y(FE_MDBN8_), 
	.A(fft_data_in[24]));
   BUFX2TS FE_MDBC7_U5210 (.Y(FE_MDBN7_), 
	.A(fft_data_in[5]));
   BUFX2TS FE_MDBC6_U5209 (.Y(FE_MDBN6_), 
	.A(fft_data_in[3]));
   BUFX2TS FE_MDBC5_U5208 (.Y(FE_MDBN5_), 
	.A(fft_data_in[2]));
   BUFX2TS FE_MDBC4_U5719 (.Y(FE_MDBN4_), 
	.A(fft_data_in[1]));
   BUFX2TS FE_MDBC3_U5677 (.Y(FE_MDBN3_), 
	.A(fft_data_in[0]));
   BUFX2TS FE_MDBC2_U5721 (.Y(FE_MDBN2_), 
	.A(fir_data_in[31]));
   BUFX2TS FE_MDBC1_U5586 (.Y(FE_MDBN1_), 
	.A(fir_data_in[29]));
   BUFX2TS FE_MDBC0_U5490 (.Y(FE_MDBN0_), 
	.A(fir_data_in[28]));
   DFFTRX1TS \mips/mips/a/accbypassA_reg  (.RN(n4444), 
	.Q(acc_bypass), 
	.D(n3440), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[31]  (.RN(n9370), 
	.Q(instruction[31]), 
	.D(\mips/mips/accfullinstruction[31] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[30]  (.RN(n9370), 
	.Q(instruction[30]), 
	.D(\mips/mips/accfullinstruction[30] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[29]  (.RN(n9370), 
	.Q(instruction[29]), 
	.D(\mips/mips/accfullinstruction[29] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[28]  (.RN(n9371), 
	.Q(instruction[28]), 
	.D(\mips/mips/accfullinstruction[28] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[27]  (.RN(n9371), 
	.Q(instruction[27]), 
	.D(\mips/mips/accfullinstruction[27] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[26]  (.RN(n9371), 
	.Q(instruction[26]), 
	.D(\mips/mips/accfullinstruction[26] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[0]  (.RN(n9371), 
	.Q(instruction[0]), 
	.D(\mips/mips/accfullinstruction[0] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[1]  (.RN(n9372), 
	.QN(n3455), 
	.Q(instruction[1]), 
	.D(\mips/mips/accfullinstruction[1] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[2]  (.RN(n9372), 
	.Q(instruction[2]), 
	.D(\mips/mips/accfullinstruction[2] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[3]  (.RN(n9372), 
	.Q(instruction[3]), 
	.D(\mips/mips/accfullinstruction[3] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[4]  (.RN(n9372), 
	.Q(instruction[4]), 
	.D(\mips/mips/accfullinstruction[4] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[5]  (.RN(n9373), 
	.Q(instruction[5]), 
	.D(\mips/mips/accfullinstruction[5] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[6]  (.RN(n9373), 
	.Q(instruction[6]), 
	.D(\mips/mips/accfullinstruction[6] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[7]  (.RN(n9373), 
	.Q(instruction[7]), 
	.D(\mips/mips/accfullinstruction[7] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[8]  (.RN(n9373), 
	.Q(instruction[8]), 
	.D(\mips/mips/accfullinstruction[8] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[9]  (.RN(n9374), 
	.Q(instruction[9]), 
	.D(\mips/mips/accfullinstruction[9] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[10]  (.RN(n9374), 
	.Q(instruction[10]), 
	.D(\mips/mips/accfullinstruction[10] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[11]  (.RN(n9374), 
	.Q(instruction[11]), 
	.D(\mips/mips/accfullinstruction[11] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[12]  (.RN(n9374), 
	.Q(instruction[12]), 
	.D(\mips/mips/accfullinstruction[12] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[13]  (.RN(n9375), 
	.Q(instruction[13]), 
	.D(\mips/mips/accfullinstruction[13] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[14]  (.RN(n9375), 
	.Q(instruction[14]), 
	.D(\mips/mips/accfullinstruction[14] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[15]  (.RN(n9375), 
	.Q(instruction[15]), 
	.D(\mips/mips/accfullinstruction[15] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[16]  (.RN(n9375), 
	.Q(instruction[16]), 
	.D(\mips/mips/accfullinstruction[16] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[17]  (.RN(n9376), 
	.Q(instruction[17]), 
	.D(\mips/mips/accfullinstruction[17] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[18]  (.RN(n9376), 
	.Q(instruction[18]), 
	.D(\mips/mips/accfullinstruction[18] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[19]  (.RN(n9376), 
	.Q(instruction[19]), 
	.D(\mips/mips/accfullinstruction[19] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[20]  (.RN(n9376), 
	.Q(instruction[20]), 
	.D(\mips/mips/accfullinstruction[20] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[21]  (.RN(n9377), 
	.Q(instruction[21]), 
	.D(\mips/mips/accfullinstruction[21] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[22]  (.RN(n9377), 
	.Q(instruction[22]), 
	.D(\mips/mips/accfullinstruction[22] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[23]  (.RN(n9377), 
	.Q(instruction[23]), 
	.D(\mips/mips/accfullinstruction[23] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[24]  (.RN(n9377), 
	.Q(instruction[24]), 
	.D(\mips/mips/accfullinstruction[24] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \mips/mips/a/fullinstructionA_reg[25]  (.RN(n9378), 
	.Q(instruction[25]), 
	.D(\mips/mips/accfullinstruction[25] ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell14/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell15/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[14] ), 
	.D(\fifo_from_fir/fifo_cell14/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell13/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell14/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[13] ), 
	.D(\fifo_from_fir/fifo_cell13/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell12/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell13/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[12] ), 
	.D(\fifo_from_fir/fifo_cell12/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell11/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell12/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[11] ), 
	.D(\fifo_from_fir/fifo_cell11/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell10/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell11/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[10] ), 
	.D(\fifo_from_fir/fifo_cell10/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell9/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell10/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[9] ), 
	.D(\fifo_from_fir/fifo_cell9/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell8/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell9/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[8] ), 
	.D(\fifo_from_fir/fifo_cell8/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell7/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell8/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[7] ), 
	.D(\fifo_from_fir/fifo_cell7/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell6/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell7/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[6] ), 
	.D(\fifo_from_fir/fifo_cell6/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell5/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell6/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[5] ), 
	.D(\fifo_from_fir/fifo_cell5/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell4/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell5/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[4] ), 
	.D(\fifo_from_fir/fifo_cell4/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell3/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell4/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[3] ), 
	.D(\fifo_from_fir/fifo_cell3/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell2/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell3/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[2] ), 
	.D(\fifo_from_fir/fifo_cell2/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell1/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell2/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[1] ), 
	.D(\fifo_from_fir/fifo_cell1/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fir/fifo_cell0/hold_token_reg  (.RN(\fifo_from_fir/fifo_cell1/data_out/N35 ), 
	.Q(\fifo_from_fir/hold[0] ), 
	.D(\fifo_from_fir/fifo_cell0/data_out/N9 ), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell1/controller/write_enable_reg  (.RN(n9542), 
	.QN(\fifo_from_fir/fifo_cell1/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell1/controller/valid_read ), 
	.D(n7598), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell2/controller/write_enable_reg  (.RN(n9542), 
	.QN(\fifo_from_fir/fifo_cell2/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell2/controller/valid_read ), 
	.D(n7593), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell3/controller/write_enable_reg  (.RN(n9543), 
	.QN(\fifo_from_fir/fifo_cell3/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell3/controller/valid_read ), 
	.D(n7588), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell4/controller/write_enable_reg  (.RN(n9545), 
	.QN(\fifo_from_fir/fifo_cell4/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell4/controller/valid_read ), 
	.D(n7583), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell5/controller/write_enable_reg  (.RN(n9543), 
	.QN(\fifo_from_fir/fifo_cell5/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell5/controller/valid_read ), 
	.D(n7578), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell6/controller/write_enable_reg  (.RN(n9545), 
	.QN(\fifo_from_fir/fifo_cell6/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell6/controller/valid_read ), 
	.D(n7573), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell7/controller/write_enable_reg  (.RN(n9544), 
	.QN(\fifo_from_fir/fifo_cell7/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell7/controller/valid_read ), 
	.D(n7568), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell8/controller/write_enable_reg  (.RN(n9544), 
	.QN(\fifo_from_fir/fifo_cell8/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell8/controller/valid_read ), 
	.D(n7563), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell9/controller/write_enable_reg  (.RN(n9544), 
	.QN(\fifo_from_fir/fifo_cell9/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell9/controller/valid_read ), 
	.D(n7558), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell10/controller/write_enable_reg  (.RN(n9543), 
	.QN(\fifo_from_fir/fifo_cell10/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell10/controller/valid_read ), 
	.D(n7553), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell11/controller/write_enable_reg  (.RN(n9543), 
	.QN(\fifo_from_fir/fifo_cell11/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell11/controller/valid_read ), 
	.D(n7548), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell12/controller/write_enable_reg  (.RN(n7618), 
	.QN(\fifo_from_fir/fifo_cell12/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell12/controller/valid_read ), 
	.D(n7543), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell13/controller/write_enable_reg  (.RN(n9547), 
	.QN(\fifo_from_fir/fifo_cell13/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell13/controller/valid_read ), 
	.D(n7538), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell14/controller/write_enable_reg  (.RN(n9538), 
	.QN(\fifo_from_fir/fifo_cell14/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell14/controller/valid_read ), 
	.D(n7533), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell15/controller/write_enable_reg  (.RN(n9539), 
	.QN(\fifo_from_fir/fifo_cell15/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell15/controller/valid_read ), 
	.D(n7528), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/addr_calc/fir_read_calc/counter/count_reg[0]  (.QN(n7955), 
	.Q(\router/addr_calc/fir_read_calc/count[0] ), 
	.E(FE_OFN1190_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N178 ), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/addr_calc/fir_write_calc/counter/count_reg[0]  (.QN(n7956), 
	.Q(\router/addr_calc/fir_write_calc/count[0] ), 
	.E(FE_OFN1179_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N178 ), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/addr_calc/fft_read_calc/counter/count_reg[0]  (.QN(n7957), 
	.Q(\router/addr_calc/fft_read_calc/count[0] ), 
	.E(FE_OFN1169_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N178 ), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/addr_calc/fft_write_calc/counter/count_reg[0]  (.QN(n7958), 
	.Q(\router/addr_calc/fft_write_calc/count[0] ), 
	.E(FE_OFN1161_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N178 ), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell0/controller/write_enable_reg  (.RN(n9537), 
	.QN(\fifo_to_fft/fifo_cell0/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell0/controller/valid_read ), 
	.D(n7231), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell15/data_out/en_reg  (.RN(n3959), 
	.Q(\fifo_to_fft/fifo_cell15/control_signal ), 
	.D(\fifo_to_fft/fifo_cell14/reg_gtok/token ), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell15/controller/write_enable_reg  (.RN(n9538), 
	.QN(\fifo_to_fft/fifo_cell15/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell15/controller/valid_read ), 
	.D(n7241), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell14/data_out/en_reg  (.RN(FE_OFN699_n3959), 
	.QN(n2891), 
	.D(\fifo_to_fft/fifo_cell13/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell14/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell15/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[14] ), 
	.D(n2891), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell14/controller/write_enable_reg  (.RN(n9537), 
	.QN(\fifo_to_fft/fifo_cell14/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell14/controller/valid_read ), 
	.D(n7246), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell13/data_out/en_reg  (.RN(FE_OFN703_n3959), 
	.QN(n2888), 
	.D(\fifo_to_fft/fifo_cell12/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell13/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell14/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[13] ), 
	.D(n2888), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell13/controller/write_enable_reg  (.RN(n9536), 
	.QN(\fifo_to_fft/fifo_cell13/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell13/controller/valid_read ), 
	.D(n7251), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell12/data_out/en_reg  (.RN(FE_OFN707_n3959), 
	.QN(n2885), 
	.D(\fifo_to_fft/fifo_cell11/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell12/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell13/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[12] ), 
	.D(n2885), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell12/controller/write_enable_reg  (.RN(n7618), 
	.QN(\fifo_to_fft/fifo_cell12/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell12/controller/valid_read ), 
	.D(n7260), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell11/data_out/en_reg  (.RN(FE_OFN707_n3959), 
	.QN(n2882), 
	.D(\fifo_to_fft/fifo_cell10/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell11/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell12/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[11] ), 
	.D(n2882), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell11/controller/write_enable_reg  (.RN(n9532), 
	.QN(\fifo_to_fft/fifo_cell11/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell11/controller/valid_read ), 
	.D(n7270), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell10/data_out/en_reg  (.RN(FE_OFN706_n3959), 
	.QN(n2879), 
	.D(\fifo_to_fft/fifo_cell9/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell10/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell11/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[10] ), 
	.D(n2879), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell10/controller/write_enable_reg  (.RN(n9532), 
	.QN(\fifo_to_fft/fifo_cell10/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell10/controller/valid_read ), 
	.D(n7275), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell9/data_out/en_reg  (.RN(FE_OFN706_n3959), 
	.QN(n2876), 
	.D(\fifo_to_fft/fifo_cell8/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell9/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell10/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[9] ), 
	.D(n2876), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell9/controller/write_enable_reg  (.RN(n9533), 
	.QN(\fifo_to_fft/fifo_cell9/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell9/controller/valid_read ), 
	.D(n7280), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell8/data_out/en_reg  (.RN(FE_OFN705_n3959), 
	.QN(n2873), 
	.D(\fifo_to_fft/fifo_cell7/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell8/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell9/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[8] ), 
	.D(n2873), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell8/controller/write_enable_reg  (.RN(n9531), 
	.QN(\fifo_to_fft/fifo_cell8/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell8/controller/valid_read ), 
	.D(n7290), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell7/data_out/en_reg  (.RN(FE_OFN708_n3959), 
	.QN(n2870), 
	.D(\fifo_to_fft/fifo_cell6/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell7/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell8/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[7] ), 
	.D(n2870), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell7/controller/write_enable_reg  (.RN(n9536), 
	.QN(\fifo_to_fft/fifo_cell7/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell7/controller/valid_read ), 
	.D(n7300), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell6/data_out/en_reg  (.RN(FE_OFN708_n3959), 
	.QN(n2867), 
	.D(\fifo_to_fft/fifo_cell5/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell6/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell7/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[6] ), 
	.D(n2867), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell6/controller/write_enable_reg  (.RN(n9532), 
	.QN(\fifo_to_fft/fifo_cell6/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell6/controller/valid_read ), 
	.D(n7305), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell5/data_out/en_reg  (.RN(FE_OFN708_n3959), 
	.QN(n2864), 
	.D(\fifo_to_fft/fifo_cell4/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell5/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell6/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[5] ), 
	.D(n2864), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell5/controller/write_enable_reg  (.RN(n9534), 
	.QN(\fifo_to_fft/fifo_cell5/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell5/controller/valid_read ), 
	.D(n7310), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell4/data_out/en_reg  (.RN(FE_OFN704_n3959), 
	.QN(n2861), 
	.D(\fifo_to_fft/fifo_cell3/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell4/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell5/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[4] ), 
	.D(n2861), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell4/controller/write_enable_reg  (.RN(n9532), 
	.QN(\fifo_to_fft/fifo_cell4/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell4/controller/valid_read ), 
	.D(n7320), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell3/data_out/en_reg  (.RN(FE_OFN704_n3959), 
	.QN(n2858), 
	.D(\fifo_to_fft/fifo_cell2/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell3/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell4/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[3] ), 
	.D(n2858), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell3/controller/write_enable_reg  (.RN(n9536), 
	.QN(\fifo_to_fft/fifo_cell3/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell3/controller/valid_read ), 
	.D(n7325), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell2/data_out/en_reg  (.RN(FE_OFN701_n3959), 
	.QN(n2855), 
	.D(\fifo_to_fft/fifo_cell1/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell2/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell3/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[2] ), 
	.D(n2855), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell2/controller/write_enable_reg  (.RN(n9535), 
	.QN(\fifo_to_fft/fifo_cell2/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell2/controller/valid_read ), 
	.D(n7330), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell1/data_out/en_reg  (.RN(FE_OFN700_n3959), 
	.QN(n2852), 
	.D(\fifo_to_fft/fifo_cell0/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fft/fifo_cell1/hold_token_reg  (.RN(\fifo_to_fft/fifo_cell2/data_out/N35 ), 
	.Q(\fifo_to_fft/hold[1] ), 
	.D(n2852), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fft/fifo_cell1/controller/write_enable_reg  (.RN(n9546), 
	.QN(\fifo_to_fft/fifo_cell1/controller/write_enable ), 
	.E(\fifo_to_fft/fifo_cell1/controller/valid_read ), 
	.D(n7340), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/data_cntl/fir_full_flag_reg  (.QN(n3470), 
	.Q(\router/data_cntl/fir_full_flag ), 
	.E(n8095), 
	.D(FE_OFN1285_router_ram_read_enable_reg), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell0/controller/write_enable_reg  (.RN(n9533), 
	.QN(\fifo_to_fir/fifo_cell0/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell0/controller/valid_read ), 
	.D(n7226), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell15/data_out/en_reg  (.RN(FE_OFN684_n4134), 
	.Q(\fifo_to_fir/fifo_cell15/control_signal ), 
	.D(\fifo_to_fir/fifo_cell14/reg_gtok/token ), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell15/controller/write_enable_reg  (.RN(n9533), 
	.QN(\fifo_to_fir/fifo_cell15/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell15/controller/valid_read ), 
	.D(n7350), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell14/data_out/en_reg  (.RN(FE_OFN695_n4134), 
	.QN(n2843), 
	.D(\fifo_to_fir/fifo_cell13/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell14/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell15/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[14] ), 
	.D(n2843), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell14/controller/write_enable_reg  (.RN(n9535), 
	.QN(\fifo_to_fir/fifo_cell14/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell14/controller/valid_read ), 
	.D(n7355), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell13/data_out/en_reg  (.RN(FE_OFN695_n4134), 
	.QN(n2840), 
	.D(\fifo_to_fir/fifo_cell12/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell13/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell14/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[13] ), 
	.D(n2840), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell13/controller/write_enable_reg  (.RN(n9533), 
	.QN(\fifo_to_fir/fifo_cell13/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell13/controller/valid_read ), 
	.D(n7360), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell12/data_out/en_reg  (.RN(FE_OFN694_n4134), 
	.QN(n2837), 
	.D(\fifo_to_fir/fifo_cell11/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell12/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell13/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[12] ), 
	.D(n2837), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell12/controller/write_enable_reg  (.RN(n9534), 
	.QN(\fifo_to_fir/fifo_cell12/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell12/controller/valid_read ), 
	.D(n7369), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell11/data_out/en_reg  (.RN(FE_OFN693_n4134), 
	.QN(n2834), 
	.D(\fifo_to_fir/fifo_cell10/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell11/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell12/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[11] ), 
	.D(n2834), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell11/controller/write_enable_reg  (.RN(n9537), 
	.QN(\fifo_to_fir/fifo_cell11/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell11/controller/valid_read ), 
	.D(n7379), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell10/data_out/en_reg  (.RN(FE_OFN693_n4134), 
	.QN(n2831), 
	.D(\fifo_to_fir/fifo_cell9/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell10/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell11/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[10] ), 
	.D(n2831), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell10/controller/write_enable_reg  (.RN(n9534), 
	.QN(\fifo_to_fir/fifo_cell10/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell10/controller/valid_read ), 
	.D(n7384), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell9/data_out/en_reg  (.RN(FE_OFN691_n4134), 
	.QN(n2828), 
	.D(\fifo_to_fir/fifo_cell8/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell9/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell10/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[9] ), 
	.D(n2828), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell9/controller/write_enable_reg  (.RN(n9534), 
	.QN(\fifo_to_fir/fifo_cell9/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell9/controller/valid_read ), 
	.D(n7389), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell8/data_out/en_reg  (.RN(FE_OFN689_n4134), 
	.QN(n2825), 
	.D(\fifo_to_fir/fifo_cell7/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell8/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell9/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[8] ), 
	.D(n2825), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell8/controller/write_enable_reg  (.RN(n9537), 
	.QN(\fifo_to_fir/fifo_cell8/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell8/controller/valid_read ), 
	.D(n7399), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell7/data_out/en_reg  (.RN(FE_OFN689_n4134), 
	.QN(n2822), 
	.D(\fifo_to_fir/fifo_cell6/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell7/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell8/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[7] ), 
	.D(n2822), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell7/controller/write_enable_reg  (.RN(n9535), 
	.QN(\fifo_to_fir/fifo_cell7/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell7/controller/valid_read ), 
	.D(n7409), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell6/data_out/en_reg  (.RN(FE_OFN688_n4134), 
	.QN(n2819), 
	.D(\fifo_to_fir/fifo_cell5/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell6/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell7/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[6] ), 
	.D(n2819), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell6/controller/write_enable_reg  (.RN(n9535), 
	.QN(\fifo_to_fir/fifo_cell6/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell6/controller/valid_read ), 
	.D(n7414), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell5/data_out/en_reg  (.RN(FE_OFN685_n4134), 
	.QN(n2816), 
	.D(\fifo_to_fir/fifo_cell4/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell5/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell6/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[5] ), 
	.D(n2816), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell5/controller/write_enable_reg  (.RN(n7618), 
	.QN(\fifo_to_fir/fifo_cell5/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell5/controller/valid_read ), 
	.D(n7419), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell4/data_out/en_reg  (.RN(FE_OFN686_n4134), 
	.QN(n2813), 
	.D(\fifo_to_fir/fifo_cell3/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell4/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell5/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[4] ), 
	.D(n2813), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell4/controller/write_enable_reg  (.RN(n9539), 
	.QN(\fifo_to_fir/fifo_cell4/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell4/controller/valid_read ), 
	.D(n7429), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell3/data_out/en_reg  (.RN(FE_OFN685_n4134), 
	.QN(n2810), 
	.D(\fifo_to_fir/fifo_cell2/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell3/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell4/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[3] ), 
	.D(n2810), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell3/controller/write_enable_reg  (.RN(n9536), 
	.QN(\fifo_to_fir/fifo_cell3/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell3/controller/valid_read ), 
	.D(n7434), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell2/data_out/en_reg  (.RN(FE_OFN684_n4134), 
	.QN(n2807), 
	.D(\fifo_to_fir/fifo_cell1/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell2/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell3/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[2] ), 
	.D(n2807), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell2/controller/write_enable_reg  (.RN(n9538), 
	.QN(\fifo_to_fir/fifo_cell2/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell2/controller/valid_read ), 
	.D(n7439), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell1/data_out/en_reg  (.RN(FE_OFN683_n4134), 
	.QN(n2804), 
	.D(\fifo_to_fir/fifo_cell0/reg_gtok/token ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_to_fir/fifo_cell1/hold_token_reg  (.RN(\fifo_to_fir/fifo_cell2/data_out/N35 ), 
	.Q(\fifo_to_fir/hold[1] ), 
	.D(n2804), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_to_fir/fifo_cell1/controller/write_enable_reg  (.RN(n9538), 
	.QN(\fifo_to_fir/fifo_cell1/controller/write_enable ), 
	.E(\fifo_to_fir/fifo_cell1/controller/valid_read ), 
	.D(n7449), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell14/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell15/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[14] ), 
	.D(\fifo_from_fft/fifo_cell14/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell13/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell14/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[13] ), 
	.D(\fifo_from_fft/fifo_cell13/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell12/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell13/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[12] ), 
	.D(\fifo_from_fft/fifo_cell12/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell11/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell12/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[11] ), 
	.D(\fifo_from_fft/fifo_cell11/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell10/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell11/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[10] ), 
	.D(\fifo_from_fft/fifo_cell10/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell9/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell10/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[9] ), 
	.D(\fifo_from_fft/fifo_cell9/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell8/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell9/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[8] ), 
	.D(\fifo_from_fft/fifo_cell8/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell7/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell8/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[7] ), 
	.D(\fifo_from_fft/fifo_cell7/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell6/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell7/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[6] ), 
	.D(\fifo_from_fft/fifo_cell6/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell5/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell6/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[5] ), 
	.D(\fifo_from_fft/fifo_cell5/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell4/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell5/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[4] ), 
	.D(\fifo_from_fft/fifo_cell4/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell3/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell4/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[3] ), 
	.D(\fifo_from_fft/fifo_cell3/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell2/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell3/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[2] ), 
	.D(\fifo_from_fft/fifo_cell2/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell1/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell2/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[1] ), 
	.D(\fifo_from_fft/fifo_cell1/data_out/N9 ), 
	.CK(clk__L1_N0));
   DFFTRX1TS \fifo_from_fft/fifo_cell0/hold_token_reg  (.RN(\fifo_from_fft/fifo_cell1/data_out/N35 ), 
	.Q(\fifo_from_fft/hold[0] ), 
	.D(\fifo_from_fft/fifo_cell0/data_out/N9 ), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell1/controller/write_enable_reg  (.RN(n9539), 
	.QN(\fifo_from_fft/fifo_cell1/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell1/controller/valid_read ), 
	.D(n7523), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell2/controller/write_enable_reg  (.RN(n9539), 
	.QN(\fifo_from_fft/fifo_cell2/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell2/controller/valid_read ), 
	.D(n7518), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell3/controller/write_enable_reg  (.RN(n9540), 
	.QN(\fifo_from_fft/fifo_cell3/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell3/controller/valid_read ), 
	.D(n7513), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell4/controller/write_enable_reg  (.RN(n9540), 
	.QN(\fifo_from_fft/fifo_cell4/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell4/controller/valid_read ), 
	.D(n7508), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell5/controller/write_enable_reg  (.RN(n9540), 
	.QN(\fifo_from_fft/fifo_cell5/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell5/controller/valid_read ), 
	.D(n7503), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell6/controller/write_enable_reg  (.RN(n9540), 
	.QN(\fifo_from_fft/fifo_cell6/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell6/controller/valid_read ), 
	.D(n7498), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell7/controller/write_enable_reg  (.RN(n9541), 
	.QN(\fifo_from_fft/fifo_cell7/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell7/controller/valid_read ), 
	.D(n7493), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell8/controller/write_enable_reg  (.RN(n9541), 
	.QN(\fifo_from_fft/fifo_cell8/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell8/controller/valid_read ), 
	.D(n7489), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell9/controller/write_enable_reg  (.RN(n9541), 
	.QN(\fifo_from_fft/fifo_cell9/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell9/controller/valid_read ), 
	.D(n7484), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell10/controller/write_enable_reg  (.RN(n9541), 
	.QN(\fifo_from_fft/fifo_cell10/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell10/controller/valid_read ), 
	.D(n7479), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell11/controller/write_enable_reg  (.RN(n9542), 
	.QN(\fifo_from_fft/fifo_cell11/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell11/controller/valid_read ), 
	.D(n7474), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell12/controller/write_enable_reg  (.RN(n9542), 
	.QN(\fifo_from_fft/fifo_cell12/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell12/controller/valid_read ), 
	.D(n7469), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell13/controller/write_enable_reg  (.RN(n9544), 
	.QN(\fifo_from_fft/fifo_cell13/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell13/controller/valid_read ), 
	.D(n7464), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell14/controller/write_enable_reg  (.RN(n9545), 
	.QN(\fifo_from_fft/fifo_cell14/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell14/controller/valid_read ), 
	.D(n7459), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell15/controller/write_enable_reg  (.RN(n9545), 
	.QN(\fifo_from_fft/fifo_cell15/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell15/controller/valid_read ), 
	.D(n7454), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/addr_calc/iir_write_calc/counter/count_reg[0]  (.QN(n7959), 
	.Q(\router/addr_calc/iir_write_calc/count[0] ), 
	.E(FE_OFN1207_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N178 ), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/addr_calc/iir_write_calc/counter/count_reg[16]  (.Q(\router/addr_calc/iir_write_calc/count[16] ), 
	.E(FE_OFN1205_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N194 ), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/addr_calc/iir_write_calc/counter/count_reg[19]  (.Q(\router/addr_calc/iir_write_calc/count[19] ), 
	.E(FE_OFN1202_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N197 ), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/addr_calc/iir_write_calc/counter/count_reg[27]  (.Q(\router/addr_calc/iir_write_calc/count[27] ), 
	.E(FE_OFN1199_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N205 ), 
	.CK(clk__L1_N0));
   EDFFX1TS \router/addr_calc/iir_write_calc/counter/count_reg[30]  (.QN(n7952), 
	.Q(\router/addr_calc/iir_write_calc/count[30] ), 
	.E(n7014), 
	.D(\router/addr_calc/iir_write_calc/counter/N208 ), 
	.CK(clk__L1_N0));
   NAND2X1TS U218 (.Y(\router/data_cntl/N138 ), 
	.B(n3469), 
	.A(n3468));
   NAND2X1TS U233 (.Y(\router/addr_calc/iir_write_calc/counter/N208 ), 
	.B(n3488), 
	.A(FE_OFN1293_iir_enable));
   NAND2X1TS U235 (.Y(\router/addr_calc/iir_write_calc/counter/N207 ), 
	.B(n3489), 
	.A(FE_OFN1295_iir_enable));
   NAND2X1TS U237 (.Y(\router/addr_calc/iir_write_calc/counter/N206 ), 
	.B(n3490), 
	.A(FE_OFN1296_iir_enable));
   NAND2X1TS U239 (.Y(\router/addr_calc/iir_write_calc/counter/N205 ), 
	.B(n3491), 
	.A(FE_OFN1296_iir_enable));
   NAND2X1TS U241 (.Y(\router/addr_calc/iir_write_calc/counter/N204 ), 
	.B(n3492), 
	.A(FE_OFN1296_iir_enable));
   NAND2X1TS U243 (.Y(\router/addr_calc/iir_write_calc/counter/N203 ), 
	.B(n3493), 
	.A(FE_OFN1293_iir_enable));
   NAND2X1TS U245 (.Y(\router/addr_calc/iir_write_calc/counter/N202 ), 
	.B(n3494), 
	.A(FE_OFN1291_iir_enable));
   NAND2X1TS U247 (.Y(\router/addr_calc/iir_write_calc/counter/N201 ), 
	.B(n3495), 
	.A(FE_OFN1291_iir_enable));
   NAND2X1TS U249 (.Y(\router/addr_calc/iir_write_calc/counter/N200 ), 
	.B(n3496), 
	.A(FE_OFN1288_iir_enable));
   NAND2X1TS U251 (.Y(\router/addr_calc/iir_write_calc/counter/N199 ), 
	.B(n3497), 
	.A(FE_OFN1290_iir_enable));
   NAND2X1TS U253 (.Y(\router/addr_calc/iir_write_calc/counter/N198 ), 
	.B(n3498), 
	.A(FE_OFN1290_iir_enable));
   NAND2X1TS U255 (.Y(\router/addr_calc/iir_write_calc/counter/N197 ), 
	.B(n3499), 
	.A(FE_OFN1292_iir_enable));
   NAND2X1TS U257 (.Y(\router/addr_calc/iir_write_calc/counter/N196 ), 
	.B(n3500), 
	.A(FE_OFN1292_iir_enable));
   NAND2X1TS U259 (.Y(\router/addr_calc/iir_write_calc/counter/N195 ), 
	.B(n3501), 
	.A(FE_OFN1292_iir_enable));
   NAND2X1TS U261 (.Y(\router/addr_calc/iir_write_calc/counter/N194 ), 
	.B(n3502), 
	.A(FE_OFN1297_iir_enable));
   NAND2X1TS U263 (.Y(\router/addr_calc/iir_write_calc/counter/N193 ), 
	.B(n3503), 
	.A(FE_OFN1294_iir_enable));
   NAND2X1TS U265 (.Y(\router/addr_calc/iir_write_calc/counter/N192 ), 
	.B(n3504), 
	.A(FE_OFN1297_iir_enable));
   NAND2X1TS U267 (.Y(\router/addr_calc/iir_write_calc/counter/N191 ), 
	.B(n3505), 
	.A(FE_OFN1297_iir_enable));
   NAND2X1TS U279 (.Y(\router/addr_calc/iir_write_calc/counter/N185 ), 
	.B(n3511), 
	.A(FE_OFN1299_iir_enable));
   NAND2X1TS U281 (.Y(\router/addr_calc/iir_write_calc/counter/N184 ), 
	.B(n3512), 
	.A(FE_OFN1299_iir_enable));
   NAND2X1TS U283 (.Y(\router/addr_calc/iir_write_calc/counter/N183 ), 
	.B(n3513), 
	.A(FE_OFN1295_iir_enable));
   NAND2X1TS U285 (.Y(\router/addr_calc/iir_write_calc/counter/N182 ), 
	.B(n3514), 
	.A(FE_OFN1295_iir_enable));
   NAND2X1TS U289 (.Y(\router/addr_calc/iir_write_calc/counter/N180 ), 
	.B(n3516), 
	.A(FE_OFN1300_iir_enable));
   NAND2X1TS U291 (.Y(\router/addr_calc/iir_write_calc/counter/N179 ), 
	.B(n3517), 
	.A(FE_OFN1300_iir_enable));
   NAND2X1TS U293 (.Y(\router/addr_calc/iir_write_calc/counter/N178 ), 
	.B(n3518), 
	.A(FE_OFN1300_iir_enable));
   NAND2X1TS U308 (.Y(\router/addr_calc/fir_write_calc/counter/N208 ), 
	.B(n3532), 
	.A(fir_enable));
   NAND2X1TS U310 (.Y(\router/addr_calc/fir_write_calc/counter/N207 ), 
	.B(n3533), 
	.A(fir_enable));
   NAND2X1TS U312 (.Y(\router/addr_calc/fir_write_calc/counter/N206 ), 
	.B(n3534), 
	.A(n9421));
   NAND2X1TS U314 (.Y(\router/addr_calc/fir_write_calc/counter/N205 ), 
	.B(n3535), 
	.A(n9421));
   NAND2X1TS U316 (.Y(\router/addr_calc/fir_write_calc/counter/N204 ), 
	.B(n3536), 
	.A(n9421));
   NAND2X1TS U318 (.Y(\router/addr_calc/fir_write_calc/counter/N203 ), 
	.B(n3537), 
	.A(n9421));
   NAND2X1TS U320 (.Y(\router/addr_calc/fir_write_calc/counter/N202 ), 
	.B(n3538), 
	.A(n9420));
   NAND2X1TS U322 (.Y(\router/addr_calc/fir_write_calc/counter/N201 ), 
	.B(n3539), 
	.A(n9420));
   NAND2X1TS U324 (.Y(\router/addr_calc/fir_write_calc/counter/N200 ), 
	.B(n3540), 
	.A(n9420));
   NAND2X1TS U326 (.Y(\router/addr_calc/fir_write_calc/counter/N199 ), 
	.B(n3541), 
	.A(n9420));
   NAND2X1TS U328 (.Y(\router/addr_calc/fir_write_calc/counter/N198 ), 
	.B(n3542), 
	.A(n9419));
   NAND2X1TS U330 (.Y(\router/addr_calc/fir_write_calc/counter/N197 ), 
	.B(n3543), 
	.A(n9419));
   NAND2X1TS U332 (.Y(\router/addr_calc/fir_write_calc/counter/N196 ), 
	.B(n3544), 
	.A(n9419));
   NAND2X1TS U334 (.Y(\router/addr_calc/fir_write_calc/counter/N195 ), 
	.B(n3545), 
	.A(n9419));
   NAND2X1TS U336 (.Y(\router/addr_calc/fir_write_calc/counter/N194 ), 
	.B(n3546), 
	.A(n9418));
   NAND2X1TS U338 (.Y(\router/addr_calc/fir_write_calc/counter/N193 ), 
	.B(n3547), 
	.A(n9418));
   NAND2X1TS U340 (.Y(\router/addr_calc/fir_write_calc/counter/N192 ), 
	.B(n3548), 
	.A(n9418));
   NAND2X1TS U342 (.Y(\router/addr_calc/fir_write_calc/counter/N191 ), 
	.B(n3549), 
	.A(n9418));
   NAND2X1TS U344 (.Y(\router/addr_calc/fir_write_calc/counter/N190 ), 
	.B(n3550), 
	.A(n9417));
   NAND2X1TS U348 (.Y(\router/addr_calc/fir_write_calc/counter/N188 ), 
	.B(n3552), 
	.A(n9417));
   NAND2X1TS U352 (.Y(\router/addr_calc/fir_write_calc/counter/N186 ), 
	.B(n3554), 
	.A(n9416));
   NAND2X1TS U354 (.Y(\router/addr_calc/fir_write_calc/counter/N185 ), 
	.B(n3555), 
	.A(n9416));
   NAND2X1TS U356 (.Y(\router/addr_calc/fir_write_calc/counter/N184 ), 
	.B(n3556), 
	.A(n9416));
   NAND2X1TS U358 (.Y(\router/addr_calc/fir_write_calc/counter/N183 ), 
	.B(n3557), 
	.A(n9416));
   NAND2X1TS U360 (.Y(\router/addr_calc/fir_write_calc/counter/N182 ), 
	.B(n3558), 
	.A(n9415));
   NAND2X1TS U362 (.Y(\router/addr_calc/fir_write_calc/counter/N181 ), 
	.B(n3559), 
	.A(n9415));
   NAND2X1TS U364 (.Y(\router/addr_calc/fir_write_calc/counter/N180 ), 
	.B(n3560), 
	.A(n9415));
   NAND2X1TS U366 (.Y(\router/addr_calc/fir_write_calc/counter/N179 ), 
	.B(n3561), 
	.A(n9415));
   NAND2X1TS U368 (.Y(\router/addr_calc/fir_write_calc/counter/N178 ), 
	.B(n3562), 
	.A(n9414));
   NAND2X1TS U381 (.Y(\router/addr_calc/fir_read_calc/counter/N209 ), 
	.B(n3573), 
	.A(n9414));
   NAND2X1TS U383 (.Y(\router/addr_calc/fir_read_calc/counter/N208 ), 
	.B(n3576), 
	.A(n9414));
   NAND2X1TS U385 (.Y(\router/addr_calc/fir_read_calc/counter/N207 ), 
	.B(n3577), 
	.A(n9414));
   NAND2X1TS U387 (.Y(\router/addr_calc/fir_read_calc/counter/N206 ), 
	.B(n3578), 
	.A(n9413));
   NAND2X1TS U389 (.Y(\router/addr_calc/fir_read_calc/counter/N205 ), 
	.B(n3579), 
	.A(n9413));
   NAND2X1TS U391 (.Y(\router/addr_calc/fir_read_calc/counter/N204 ), 
	.B(n3580), 
	.A(n9413));
   NAND2X1TS U393 (.Y(\router/addr_calc/fir_read_calc/counter/N203 ), 
	.B(n3581), 
	.A(n9412));
   NAND2X1TS U395 (.Y(\router/addr_calc/fir_read_calc/counter/N202 ), 
	.B(n3582), 
	.A(n9412));
   NAND2X1TS U397 (.Y(\router/addr_calc/fir_read_calc/counter/N201 ), 
	.B(n3583), 
	.A(n9412));
   NAND2X1TS U399 (.Y(\router/addr_calc/fir_read_calc/counter/N200 ), 
	.B(n3584), 
	.A(n9412));
   NAND2X1TS U401 (.Y(\router/addr_calc/fir_read_calc/counter/N199 ), 
	.B(n3585), 
	.A(n9411));
   NAND2X1TS U403 (.Y(\router/addr_calc/fir_read_calc/counter/N198 ), 
	.B(n3586), 
	.A(n9411));
   NAND2X1TS U405 (.Y(\router/addr_calc/fir_read_calc/counter/N197 ), 
	.B(n3587), 
	.A(n9411));
   NAND2X1TS U407 (.Y(\router/addr_calc/fir_read_calc/counter/N196 ), 
	.B(n3588), 
	.A(n9411));
   NAND2X1TS U409 (.Y(\router/addr_calc/fir_read_calc/counter/N195 ), 
	.B(n3589), 
	.A(n9615));
   NAND2X1TS U411 (.Y(\router/addr_calc/fir_read_calc/counter/N194 ), 
	.B(n3590), 
	.A(fir_enable));
   NAND2X1TS U413 (.Y(\router/addr_calc/fir_read_calc/counter/N193 ), 
	.B(n3591), 
	.A(fir_enable));
   NAND2X1TS U415 (.Y(\router/addr_calc/fir_read_calc/counter/N192 ), 
	.B(n3592), 
	.A(n9615));
   NAND2X1TS U417 (.Y(\router/addr_calc/fir_read_calc/counter/N191 ), 
	.B(n3593), 
	.A(n9410));
   NAND2X1TS U419 (.Y(\router/addr_calc/fir_read_calc/counter/N190 ), 
	.B(n3594), 
	.A(n9410));
   NAND2X1TS U423 (.Y(\router/addr_calc/fir_read_calc/counter/N188 ), 
	.B(n3596), 
	.A(n9410));
   NAND2X1TS U427 (.Y(\router/addr_calc/fir_read_calc/counter/N186 ), 
	.B(n3598), 
	.A(n9409));
   NAND2X1TS U429 (.Y(\router/addr_calc/fir_read_calc/counter/N185 ), 
	.B(n3599), 
	.A(n9409));
   NAND2X1TS U431 (.Y(\router/addr_calc/fir_read_calc/counter/N184 ), 
	.B(n3600), 
	.A(n9409));
   NAND2X1TS U433 (.Y(\router/addr_calc/fir_read_calc/counter/N183 ), 
	.B(n3601), 
	.A(n9409));
   NAND2X1TS U435 (.Y(\router/addr_calc/fir_read_calc/counter/N182 ), 
	.B(n3602), 
	.A(n9408));
   NAND2X1TS U437 (.Y(\router/addr_calc/fir_read_calc/counter/N181 ), 
	.B(n3603), 
	.A(n9408));
   NAND2X1TS U439 (.Y(\router/addr_calc/fir_read_calc/counter/N180 ), 
	.B(n3604), 
	.A(n9408));
   NAND2X1TS U441 (.Y(\router/addr_calc/fir_read_calc/counter/N179 ), 
	.B(n3605), 
	.A(n9408));
   NAND2X1TS U456 (.Y(\router/addr_calc/fft_write_calc/counter/N209 ), 
	.B(n3617), 
	.A(n9449));
   NAND2X1TS U458 (.Y(\router/addr_calc/fft_write_calc/counter/N208 ), 
	.B(n3620), 
	.A(fft_enable));
   NAND2X1TS U460 (.Y(\router/addr_calc/fft_write_calc/counter/N207 ), 
	.B(n3621), 
	.A(n9449));
   NAND2X1TS U462 (.Y(\router/addr_calc/fft_write_calc/counter/N206 ), 
	.B(n3622), 
	.A(n9448));
   NAND2X1TS U464 (.Y(\router/addr_calc/fft_write_calc/counter/N205 ), 
	.B(n3623), 
	.A(n9449));
   NAND2X1TS U466 (.Y(\router/addr_calc/fft_write_calc/counter/N204 ), 
	.B(n3624), 
	.A(n9449));
   NAND2X1TS U468 (.Y(\router/addr_calc/fft_write_calc/counter/N203 ), 
	.B(n3625), 
	.A(n9448));
   NAND2X1TS U470 (.Y(\router/addr_calc/fft_write_calc/counter/N202 ), 
	.B(n3626), 
	.A(n9448));
   NAND2X1TS U472 (.Y(\router/addr_calc/fft_write_calc/counter/N201 ), 
	.B(n3627), 
	.A(n9448));
   NAND2X1TS U474 (.Y(\router/addr_calc/fft_write_calc/counter/N200 ), 
	.B(n3628), 
	.A(n9447));
   NAND2X1TS U476 (.Y(\router/addr_calc/fft_write_calc/counter/N199 ), 
	.B(n3629), 
	.A(n9447));
   NAND2X1TS U478 (.Y(\router/addr_calc/fft_write_calc/counter/N198 ), 
	.B(n3630), 
	.A(n9447));
   NAND2X1TS U480 (.Y(\router/addr_calc/fft_write_calc/counter/N197 ), 
	.B(n3631), 
	.A(n9446));
   NAND2X1TS U482 (.Y(\router/addr_calc/fft_write_calc/counter/N196 ), 
	.B(n3632), 
	.A(n9447));
   NAND2X1TS U484 (.Y(\router/addr_calc/fft_write_calc/counter/N195 ), 
	.B(n3633), 
	.A(n9446));
   NAND2X1TS U486 (.Y(\router/addr_calc/fft_write_calc/counter/N194 ), 
	.B(n3634), 
	.A(n9445));
   NAND2X1TS U488 (.Y(\router/addr_calc/fft_write_calc/counter/N193 ), 
	.B(n3635), 
	.A(n9446));
   NAND2X1TS U490 (.Y(\router/addr_calc/fft_write_calc/counter/N192 ), 
	.B(n3636), 
	.A(n9446));
   NAND2X1TS U492 (.Y(\router/addr_calc/fft_write_calc/counter/N191 ), 
	.B(n3637), 
	.A(n9445));
   NAND2X1TS U494 (.Y(\router/addr_calc/fft_write_calc/counter/N190 ), 
	.B(n3638), 
	.A(n9445));
   NAND2X1TS U498 (.Y(\router/addr_calc/fft_write_calc/counter/N188 ), 
	.B(n3640), 
	.A(n9444));
   NAND2X1TS U502 (.Y(\router/addr_calc/fft_write_calc/counter/N186 ), 
	.B(n3642), 
	.A(n9444));
   NAND2X1TS U504 (.Y(\router/addr_calc/fft_write_calc/counter/N185 ), 
	.B(n3643), 
	.A(n9444));
   NAND2X1TS U506 (.Y(\router/addr_calc/fft_write_calc/counter/N184 ), 
	.B(n3644), 
	.A(n9443));
   NAND2X1TS U508 (.Y(\router/addr_calc/fft_write_calc/counter/N183 ), 
	.B(n3645), 
	.A(n9443));
   NAND2X1TS U510 (.Y(\router/addr_calc/fft_write_calc/counter/N182 ), 
	.B(n3646), 
	.A(n9443));
   NAND2X1TS U512 (.Y(\router/addr_calc/fft_write_calc/counter/N181 ), 
	.B(n3647), 
	.A(n9443));
   NAND2X1TS U514 (.Y(\router/addr_calc/fft_write_calc/counter/N180 ), 
	.B(n3648), 
	.A(n9442));
   NAND2X1TS U516 (.Y(\router/addr_calc/fft_write_calc/counter/N179 ), 
	.B(n3649), 
	.A(n9442));
   NAND2X1TS U518 (.Y(\router/addr_calc/fft_write_calc/counter/N178 ), 
	.B(n3650), 
	.A(n9442));
   NAND2X1TS U531 (.Y(\router/addr_calc/fft_read_calc/counter/N209 ), 
	.B(n3661), 
	.A(n9442));
   NAND2X1TS U533 (.Y(\router/addr_calc/fft_read_calc/counter/N208 ), 
	.B(n3664), 
	.A(n9441));
   NAND2X1TS U535 (.Y(\router/addr_calc/fft_read_calc/counter/N207 ), 
	.B(n3665), 
	.A(n9441));
   NAND2X1TS U537 (.Y(\router/addr_calc/fft_read_calc/counter/N206 ), 
	.B(n3666), 
	.A(n9441));
   NAND2X1TS U539 (.Y(\router/addr_calc/fft_read_calc/counter/N205 ), 
	.B(n3667), 
	.A(n9440));
   NAND2X1TS U541 (.Y(\router/addr_calc/fft_read_calc/counter/N204 ), 
	.B(n3668), 
	.A(n9440));
   NAND2X1TS U543 (.Y(\router/addr_calc/fft_read_calc/counter/N203 ), 
	.B(n3669), 
	.A(n9440));
   NAND2X1TS U545 (.Y(\router/addr_calc/fft_read_calc/counter/N202 ), 
	.B(n3670), 
	.A(n9440));
   NAND2X1TS U547 (.Y(\router/addr_calc/fft_read_calc/counter/N201 ), 
	.B(n3671), 
	.A(n9439));
   NAND2X1TS U551 (.Y(\router/addr_calc/fft_read_calc/counter/N199 ), 
	.B(n3673), 
	.A(n9439));
   NAND2X1TS U555 (.Y(\router/addr_calc/fft_read_calc/counter/N197 ), 
	.B(n3675), 
	.A(n9438));
   NAND2X1TS U557 (.Y(\router/addr_calc/fft_read_calc/counter/N196 ), 
	.B(n3676), 
	.A(n9438));
   NAND2X1TS U559 (.Y(\router/addr_calc/fft_read_calc/counter/N195 ), 
	.B(n3677), 
	.A(n9438));
   NAND2X1TS U561 (.Y(\router/addr_calc/fft_read_calc/counter/N194 ), 
	.B(n3678), 
	.A(n9438));
   NAND2X1TS U563 (.Y(\router/addr_calc/fft_read_calc/counter/N193 ), 
	.B(n3679), 
	.A(n9437));
   NAND2X1TS U565 (.Y(\router/addr_calc/fft_read_calc/counter/N192 ), 
	.B(n3680), 
	.A(n9437));
   NAND2X1TS U567 (.Y(\router/addr_calc/fft_read_calc/counter/N191 ), 
	.B(n3681), 
	.A(n9437));
   NAND2X1TS U569 (.Y(\router/addr_calc/fft_read_calc/counter/N190 ), 
	.B(n3682), 
	.A(n9437));
   NAND2X1TS U573 (.Y(\router/addr_calc/fft_read_calc/counter/N188 ), 
	.B(n3684), 
	.A(n9436));
   NAND2X1TS U577 (.Y(\router/addr_calc/fft_read_calc/counter/N186 ), 
	.B(n3686), 
	.A(n9441));
   NAND2X1TS U579 (.Y(\router/addr_calc/fft_read_calc/counter/N185 ), 
	.B(n3687), 
	.A(n9436));
   NAND2X1TS U581 (.Y(\router/addr_calc/fft_read_calc/counter/N184 ), 
	.B(n3688), 
	.A(fft_enable));
   NAND2X1TS U583 (.Y(\router/addr_calc/fft_read_calc/counter/N183 ), 
	.B(n3689), 
	.A(fft_enable));
   NAND2X1TS U585 (.Y(\router/addr_calc/fft_read_calc/counter/N182 ), 
	.B(n3690), 
	.A(fft_enable));
   NAND2X1TS U587 (.Y(\router/addr_calc/fft_read_calc/counter/N181 ), 
	.B(n3691), 
	.A(n9614));
   NAND2X1TS U589 (.Y(\router/addr_calc/fft_read_calc/counter/N180 ), 
	.B(n3692), 
	.A(n9435));
   NAND2X1TS U591 (.Y(\router/addr_calc/fft_read_calc/counter/N179 ), 
	.B(n3693), 
	.A(n9435));
   NAND2X1TS U593 (.Y(\router/addr_calc/fft_read_calc/counter/N178 ), 
	.B(n3694), 
	.A(n9435));
   AOI222XLTS U656 (.Y(n3742), 
	.C1(fir_data_in[11]), 
	.C0(FE_OFN754_n3722), 
	.B1(fft_data_in[11]), 
	.B0(FE_OFN764_n3721), 
	.A1(\router/data_cntl/data_in[11] ), 
	.A0(FE_OFN775_n3720));
   AOI222XLTS U658 (.Y(n3743), 
	.C1(fir_data_in[10]), 
	.C0(FE_OFN754_n3722), 
	.B1(fft_data_in[10]), 
	.B0(FE_OFN764_n3721), 
	.A1(\router/data_cntl/data_in[10] ), 
	.A0(FE_OFN775_n3720));
   AOI222XLTS U670 (.Y(n3749), 
	.C1(fir_data_in[4]), 
	.C0(FE_OFN748_n3722), 
	.B1(fft_data_in[4]), 
	.B0(FE_OFN758_n3721), 
	.A1(\router/data_cntl/data_in[4] ), 
	.A0(FE_OFN769_n3720));
   NOR3BX1TS U688 (.Y(n3763), 
	.C(n3772), 
	.B(\fifo_from_fir/tok_xnor_put ), 
	.AN(\fifo_from_fir/fifo_cell0/reg_ptok/N29 ));
   NOR3BX1TS U734 (.Y(n3783), 
	.C(n3792), 
	.B(\fifo_from_fft/tok_xnor_put ), 
	.AN(\fifo_from_fft/fifo_cell0/reg_ptok/N29 ));
   NOR3BX1TS U929 (.Y(n3814), 
	.C(n4006), 
	.B(\fifo_to_fft/tok_xnor_put ), 
	.AN(\fifo_to_fft/fifo_cell0/reg_ptok/N29 ));
   AOI21X1TS U950 (.Y(n4023), 
	.B0(n4004), 
	.A1(\fifo_to_fft/fifo_cell0/reg_ptok/N29 ), 
	.A0(FE_OFN729_n8058));
   NOR3BX1TS U1073 (.Y(n3803), 
	.C(n4181), 
	.B(\fifo_to_fir/tok_xnor_put ), 
	.AN(\fifo_to_fir/fifo_cell0/reg_ptok/N29 ));
   AOI21X1TS U1094 (.Y(n4198), 
	.B0(n4179), 
	.A1(\fifo_to_fir/fifo_cell0/reg_ptok/N29 ), 
	.A0(FE_OFN732_n8057));
   NOR4XLTS U1105 (.Y(n4202), 
	.D(FE_OFN985_n9431), 
	.C(n4204), 
	.B(n4203), 
	.A(FE_OFN843_n7619));
   AO22X1TS U1499 (.Y(n5757), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[13] ), 
	.B0(FE_OFN159_n4496), 
	.A1(FE_OFN1550_acc_fft_data_in_13_), 
	.A0(FE_OFN167_n4495));
   AO22X1TS U1867 (.Y(n6095), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[15] ), 
	.B0(FE_OFN293_n4556), 
	.A1(FE_OFN1538_acc_fft_data_in_15_), 
	.A0(FE_OFN311_n4555));
   AOI21X1TS U2017 (.Y(n4595), 
	.B0(n3789), 
	.A1(\fifo_from_fft/fifo_cell0/reg_ptok/N29 ), 
	.A0(FE_OFN696_n8052));
   AO22X1TS U2130 (.Y(n6286), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[13] ), 
	.B0(FE_OFN495_n4682), 
	.A1(FE_OFN1731_acc_fir_data_in_13_), 
	.A0(FE_OFN507_n4681));
   AO22X1TS U2498 (.Y(n6624), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[15] ), 
	.B0(FE_OFN639_n4742), 
	.A1(FE_OFN1723_acc_fir_data_in_15_), 
	.A0(FE_OFN651_n4741));
   AOI21X1TS U2648 (.Y(n4781), 
	.B0(n3769), 
	.A1(\fifo_from_fir/fifo_cell0/reg_ptok/N29 ), 
	.A0(FE_OFN681_n8050));
   NAND2X1TS U2720 (.Y(n3838), 
	.B(n3835), 
	.A(n3834));
   OAI33XLTS U2730 (.Y(n6764), 
	.B2(\router/iir_write_done ), 
	.B1(n4456), 
	.B0(FE_OFN839_n7619), 
	.A2(n4449), 
	.A1(n4457), 
	.A0(n9390));
   NAND2X1TS U2734 (.Y(n4457), 
	.B(n4200), 
	.A(n3846));
   NAND2X1TS U2735 (.Y(n4200), 
	.B(n4841), 
	.A(instruction[1]));
   NAND2X1TS U3387 (.Y(n5207), 
	.B(n4132), 
	.A(\fifo_to_fir/fifo_cell1/data_out/N35 ));
   XNOR2X1TS U3400 (.Y(n5213), 
	.B(n5215), 
	.A(n5214));
   XOR2X1TS U3401 (.Y(n5215), 
	.B(n5217), 
	.A(n5216));
   XNOR2X1TS U3402 (.Y(n5217), 
	.B(n5218), 
	.A(n4123));
   XOR2X1TS U3408 (.Y(n5216), 
	.B(n5220), 
	.A(n5219));
   NAND2X1TS U3413 (.Y(n4113), 
	.B(FE_OFN686_n4134), 
	.A(\fifo_to_fir/fifo_cell3/reg_gtok/token ));
   XOR2X1TS U3419 (.Y(n5214), 
	.B(n5222), 
	.A(n5221));
   XOR2X1TS U3420 (.Y(n5222), 
	.B(n5224), 
	.A(n5223));
   XOR2X1TS U3431 (.Y(n5221), 
	.B(n5226), 
	.A(n5225));
   NAND2X1TS U3530 (.Y(n5249), 
	.B(n3957), 
	.A(\fifo_to_fft/fifo_cell1/data_out/N35 ));
   XNOR2X1TS U3544 (.Y(n5255), 
	.B(n5257), 
	.A(n5256));
   XOR2X1TS U3545 (.Y(n5257), 
	.B(n5259), 
	.A(n5258));
   XNOR2X1TS U3546 (.Y(n5259), 
	.B(n5260), 
	.A(n3948));
   XOR2X1TS U3552 (.Y(n5258), 
	.B(n5262), 
	.A(n5261));
   XOR2X1TS U3563 (.Y(n5256), 
	.B(n5264), 
	.A(n5263));
   XOR2X1TS U3564 (.Y(n5264), 
	.B(n5266), 
	.A(n5265));
   XOR2X1TS U3575 (.Y(n5263), 
	.B(n5268), 
	.A(n5267));
   NOR2X1TS U3673 (.Y(n4759), 
	.B(n5288), 
	.A(n8877));
   NOR2X1TS U3816 (.Y(n4573), 
	.B(n5327), 
	.A(n8844));
   TLATXLTS \mips/mips/a/countflag_reg  (.QN(n3440), 
	.Q(\mips/mips/a/countflag ), 
	.G(\mips/mips/a/N50 ), 
	.D(\mips/mips/a/N49 ));
   TLATXLTS \router/data_cntl/data_from_iir_reg  (.QN(n2634), 
	.Q(\router/data_from_iir ), 
	.G(\router/data_cntl/N142 ), 
	.D(n7606));
   TLATXLTS \router/data_cntl/data_to_fir_reg  (.QN(n3843), 
	.Q(\router/data_to_fir ), 
	.G(\router/data_cntl/N138 ), 
	.D(\router/data_cntl/N137 ));
   TLATXLTS \router/data_cntl/data_from_fft_reg  (.QN(n3840), 
	.Q(\router/data_from_fft ), 
	.G(\router/data_cntl/N134 ), 
	.D(\router/data_cntl/N133 ));
   TLATXLTS \router/data_cntl/data_to_fft_reg  (.QN(n3841), 
	.Q(\router/data_to_fft ), 
	.G(\router/data_cntl/N134 ), 
	.D(\router/data_cntl/N135 ));
   TLATXLTS \router/data_cntl/data_from_fir_reg  (.QN(n2633), 
	.Q(\router/data_from_fir ), 
	.G(\router/data_cntl/N138 ), 
	.D(\router/data_cntl/N139 ));
   DFFQX1TS \fifo_to_fft/fifo_cell0/data_out/en_reg  (.Q(\fifo_to_fft/fifo_cell0/control_signal ), 
	.D(\fifo_to_fft/fifo_cell0/data_out/N35 ), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell0/data_out/en_reg  (.Q(\fifo_to_fir/fifo_cell0/control_signal ), 
	.D(\fifo_to_fir/fifo_cell0/data_out/N35 ), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell0/hold_token_reg  (.Q(\fifo_to_fir/hold[0] ), 
	.D(\fifo_to_fir/fifo_cell0/N7 ), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell0/hold_token_reg  (.Q(\fifo_to_fft/hold[0] ), 
	.D(\fifo_to_fft/fifo_cell0/N7 ), 
	.CK(clk__L1_N0));
   DFFQX1TS \mips/mips/a/count_reg[0]  (.Q(\mips/mips/a/count[0] ), 
	.D(n5701), 
	.CK(clk__L1_N0));
   DFFXLTS \mips/mips/a/count_reg[1]  (.QN(n4441), 
	.D(n5700), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell0/reg_ptok/out_valid_get_reg  (.RN(n5288), 
	.QN(\fifo_from_fir/fifo_cell0/reg_ptok/out_valid_get ), 
	.D(n9547), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell0/reg_ptok/out_valid_get_reg  (.RN(n5208), 
	.QN(\fifo_to_fir/fifo_cell0/reg_ptok/out_valid_get ), 
	.D(n9547), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell0/reg_ptok/out_valid_get_reg  (.RN(n5327), 
	.QN(\fifo_from_fft/fifo_cell0/reg_ptok/out_valid_get ), 
	.D(n9546), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell0/reg_ptok/out_valid_get_reg  (.RN(n5250), 
	.QN(\fifo_to_fft/fifo_cell0/reg_ptok/out_valid_get ), 
	.D(n9547), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[31] ), 
	.D(n5385), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[30] ), 
	.D(n5386), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[29] ), 
	.D(n5387), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[28] ), 
	.D(n5388), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[27] ), 
	.D(n5389), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[26] ), 
	.D(n5390), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[25] ), 
	.D(n5391), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[24] ), 
	.D(n5392), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[23] ), 
	.D(n5393), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[22] ), 
	.D(n5394), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[21] ), 
	.D(n5395), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[20] ), 
	.D(n5396), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[19] ), 
	.D(n5397), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[18] ), 
	.D(n5398), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[17] ), 
	.D(n5399), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[16] ), 
	.D(n5400), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[15] ), 
	.D(n5401), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[14] ), 
	.D(n5402), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[13] ), 
	.D(n5403), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[12] ), 
	.D(n5404), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[11] ), 
	.D(n5405), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[10] ), 
	.D(n5406), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[9] ), 
	.D(n5407), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[8] ), 
	.D(n5408), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[7] ), 
	.D(n5409), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[6] ), 
	.D(n5410), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[5] ), 
	.D(n5411), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[4] ), 
	.D(n5412), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[3] ), 
	.D(n5413), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[2] ), 
	.D(n5414), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[1] ), 
	.D(n5415), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell0/sr_out[0] ), 
	.D(n5416), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[31] ), 
	.D(n6710), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[30] ), 
	.D(n6711), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[29] ), 
	.D(n6712), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[28] ), 
	.D(n6713), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[27] ), 
	.D(n6714), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[26] ), 
	.D(n6715), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[25] ), 
	.D(n6716), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[24] ), 
	.D(n6717), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[23] ), 
	.D(n6718), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[22] ), 
	.D(n6719), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[21] ), 
	.D(n6720), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[20] ), 
	.D(n6721), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[19] ), 
	.D(n6722), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[18] ), 
	.D(n6723), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[17] ), 
	.D(n6724), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[16] ), 
	.D(n6725), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[15] ), 
	.D(n6726), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[14] ), 
	.D(n6727), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[13] ), 
	.D(n6728), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[12] ), 
	.D(n6729), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[11] ), 
	.D(n6730), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[10] ), 
	.D(n6731), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[9] ), 
	.D(n6732), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[8] ), 
	.D(n6733), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[7] ), 
	.D(n6734), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[6] ), 
	.D(n6735), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[5] ), 
	.D(n6736), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[4] ), 
	.D(n6737), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[3] ), 
	.D(n6738), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[2] ), 
	.D(n6739), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[1] ), 
	.D(n6740), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell1/sr_out[0] ), 
	.D(n6741), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[31] ), 
	.D(n6676), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[30] ), 
	.D(n6677), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[29] ), 
	.D(n6678), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[28] ), 
	.D(n6679), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[27] ), 
	.D(n6680), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[26] ), 
	.D(n6681), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[25] ), 
	.D(n6682), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[24] ), 
	.D(n6683), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[23] ), 
	.D(n6684), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[22] ), 
	.D(n6685), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[21] ), 
	.D(n6686), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[20] ), 
	.D(n6687), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[19] ), 
	.D(n6688), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[18] ), 
	.D(n6689), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[17] ), 
	.D(n6690), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[16] ), 
	.D(n6691), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[15] ), 
	.D(n6692), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[14] ), 
	.D(n6693), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[13] ), 
	.D(n6694), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[12] ), 
	.D(n6695), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[11] ), 
	.D(n6696), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[10] ), 
	.D(n6697), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[9] ), 
	.D(n6698), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[8] ), 
	.D(n6699), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[7] ), 
	.D(n6700), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[6] ), 
	.D(n6701), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[5] ), 
	.D(n6702), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[4] ), 
	.D(n6703), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[3] ), 
	.D(n6704), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[2] ), 
	.D(n6705), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[1] ), 
	.D(n6706), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell2/sr_out[0] ), 
	.D(n6707), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[31] ), 
	.D(n6642), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[30] ), 
	.D(n6643), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[29] ), 
	.D(n6644), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[28] ), 
	.D(n6645), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[27] ), 
	.D(n6646), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[26] ), 
	.D(n6647), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[25] ), 
	.D(n6648), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[24] ), 
	.D(n6649), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[23] ), 
	.D(n6650), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[22] ), 
	.D(n6651), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[21] ), 
	.D(n6652), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[20] ), 
	.D(n6653), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[19] ), 
	.D(n6654), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[18] ), 
	.D(n6655), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[17] ), 
	.D(n6656), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[16] ), 
	.D(n6657), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[15] ), 
	.D(n6658), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[14] ), 
	.D(n6659), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[13] ), 
	.D(n6660), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[12] ), 
	.D(n6661), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[11] ), 
	.D(n6662), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[10] ), 
	.D(n6663), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[9] ), 
	.D(n6664), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[8] ), 
	.D(n6665), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[7] ), 
	.D(n6666), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[6] ), 
	.D(n6667), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[5] ), 
	.D(n6668), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[4] ), 
	.D(n6669), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[3] ), 
	.D(n6670), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[2] ), 
	.D(n6671), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[1] ), 
	.D(n6672), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell3/sr_out[0] ), 
	.D(n6673), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[31] ), 
	.D(n6608), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[30] ), 
	.D(n6609), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[29] ), 
	.D(n6610), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[28] ), 
	.D(n6611), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[27] ), 
	.D(n6612), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[26] ), 
	.D(n6613), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[25] ), 
	.D(n6614), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[24] ), 
	.D(n6615), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[23] ), 
	.D(n6616), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[22] ), 
	.D(n6617), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[21] ), 
	.D(n6618), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[20] ), 
	.D(n6619), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[19] ), 
	.D(n6620), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[18] ), 
	.D(n6621), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[17] ), 
	.D(n6622), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[16] ), 
	.D(n6623), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[15] ), 
	.D(n6624), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[14] ), 
	.D(n6625), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[13] ), 
	.D(n6626), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[12] ), 
	.D(n6627), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[11] ), 
	.D(n6628), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[10] ), 
	.D(n6629), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[9] ), 
	.D(n6630), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[8] ), 
	.D(n6631), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[7] ), 
	.D(n6632), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[6] ), 
	.D(n6633), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[5] ), 
	.D(n6634), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[4] ), 
	.D(n6635), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[3] ), 
	.D(n6636), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[2] ), 
	.D(n6637), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[1] ), 
	.D(n6638), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell4/sr_out[0] ), 
	.D(n6639), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[31] ), 
	.D(n6574), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[30] ), 
	.D(n6575), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[29] ), 
	.D(n6576), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[28] ), 
	.D(n6577), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[27] ), 
	.D(n6578), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[26] ), 
	.D(n6579), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[25] ), 
	.D(n6580), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[24] ), 
	.D(n6581), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[23] ), 
	.D(n6582), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[22] ), 
	.D(n6583), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[21] ), 
	.D(n6584), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[20] ), 
	.D(n6585), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[19] ), 
	.D(n6586), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[18] ), 
	.D(n6587), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[17] ), 
	.D(n6588), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[16] ), 
	.D(n6589), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[15] ), 
	.D(n6590), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[14] ), 
	.D(n6591), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[13] ), 
	.D(n6592), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[12] ), 
	.D(n6593), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[11] ), 
	.D(n6594), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[10] ), 
	.D(n6595), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[9] ), 
	.D(n6596), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[8] ), 
	.D(n6597), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[7] ), 
	.D(n6598), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[6] ), 
	.D(n6599), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[5] ), 
	.D(n6600), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[4] ), 
	.D(n6601), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[3] ), 
	.D(n6602), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[2] ), 
	.D(n6603), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[1] ), 
	.D(n6604), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell5/sr_out[0] ), 
	.D(n6605), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[31] ), 
	.D(n6540), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[30] ), 
	.D(n6541), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[29] ), 
	.D(n6542), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[28] ), 
	.D(n6543), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[27] ), 
	.D(n6544), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[26] ), 
	.D(n6545), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[25] ), 
	.D(n6546), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[24] ), 
	.D(n6547), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[23] ), 
	.D(n6548), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[22] ), 
	.D(n6549), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[21] ), 
	.D(n6550), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[20] ), 
	.D(n6551), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[19] ), 
	.D(n6552), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[18] ), 
	.D(n6553), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[17] ), 
	.D(n6554), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[16] ), 
	.D(n6555), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[15] ), 
	.D(n6556), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[14] ), 
	.D(n6557), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[13] ), 
	.D(n6558), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[12] ), 
	.D(n6559), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[11] ), 
	.D(n6560), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[10] ), 
	.D(n6561), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[9] ), 
	.D(n6562), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[8] ), 
	.D(n6563), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[7] ), 
	.D(n6564), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[6] ), 
	.D(n6565), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[5] ), 
	.D(n6566), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[4] ), 
	.D(n6567), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[3] ), 
	.D(n6568), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[2] ), 
	.D(n6569), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[1] ), 
	.D(n6570), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell6/sr_out[0] ), 
	.D(n6571), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[31] ), 
	.D(n6506), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[30] ), 
	.D(n6507), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[29] ), 
	.D(n6508), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[28] ), 
	.D(n6509), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[27] ), 
	.D(n6510), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[26] ), 
	.D(n6511), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[25] ), 
	.D(n6512), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[24] ), 
	.D(n6513), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[23] ), 
	.D(n6514), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[22] ), 
	.D(n6515), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[21] ), 
	.D(n6516), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[20] ), 
	.D(n6517), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[19] ), 
	.D(n6518), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[18] ), 
	.D(n6519), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[17] ), 
	.D(n6520), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[16] ), 
	.D(n6521), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[15] ), 
	.D(n6522), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[14] ), 
	.D(n6523), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[13] ), 
	.D(n6524), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[12] ), 
	.D(n6525), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[11] ), 
	.D(n6526), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[10] ), 
	.D(n6527), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[9] ), 
	.D(n6528), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[8] ), 
	.D(n6529), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[7] ), 
	.D(n6530), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[6] ), 
	.D(n6531), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[5] ), 
	.D(n6532), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[4] ), 
	.D(n6533), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[3] ), 
	.D(n6534), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[2] ), 
	.D(n6535), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[1] ), 
	.D(n6536), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell7/sr_out[0] ), 
	.D(n6537), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[31] ), 
	.D(n6472), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[30] ), 
	.D(n6473), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[29] ), 
	.D(n6474), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[28] ), 
	.D(n6475), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[27] ), 
	.D(n6476), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[26] ), 
	.D(n6477), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[25] ), 
	.D(n6478), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[24] ), 
	.D(n6479), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[23] ), 
	.D(n6480), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[22] ), 
	.D(n6481), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[21] ), 
	.D(n6482), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[20] ), 
	.D(n6483), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[19] ), 
	.D(n6484), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[18] ), 
	.D(n6485), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[17] ), 
	.D(n6486), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[16] ), 
	.D(n6487), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[15] ), 
	.D(n6488), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[14] ), 
	.D(n6489), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[13] ), 
	.D(n6490), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[12] ), 
	.D(n6491), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[11] ), 
	.D(n6492), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[10] ), 
	.D(n6493), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[9] ), 
	.D(n6494), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[8] ), 
	.D(n6495), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[7] ), 
	.D(n6496), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[6] ), 
	.D(n6497), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[5] ), 
	.D(n6498), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[4] ), 
	.D(n6499), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[3] ), 
	.D(n6500), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[2] ), 
	.D(n6501), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[1] ), 
	.D(n6502), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell8/sr_out[0] ), 
	.D(n6503), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[31] ), 
	.D(n6438), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[30] ), 
	.D(n6439), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[29] ), 
	.D(n6440), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[28] ), 
	.D(n6441), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[27] ), 
	.D(n6442), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[26] ), 
	.D(n6443), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[25] ), 
	.D(n6444), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[24] ), 
	.D(n6445), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[23] ), 
	.D(n6446), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[22] ), 
	.D(n6447), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[21] ), 
	.D(n6448), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[20] ), 
	.D(n6449), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[19] ), 
	.D(n6450), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[18] ), 
	.D(n6451), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[17] ), 
	.D(n6452), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[16] ), 
	.D(n6453), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[15] ), 
	.D(n6454), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[14] ), 
	.D(n6455), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[13] ), 
	.D(n6456), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[12] ), 
	.D(n6457), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[11] ), 
	.D(n6458), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[10] ), 
	.D(n6459), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[9] ), 
	.D(n6460), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[8] ), 
	.D(n6461), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[7] ), 
	.D(n6462), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[6] ), 
	.D(n6463), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[5] ), 
	.D(n6464), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[4] ), 
	.D(n6465), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[3] ), 
	.D(n6466), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[2] ), 
	.D(n6467), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[1] ), 
	.D(n6468), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell9/sr_out[0] ), 
	.D(n6469), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[31] ), 
	.D(n6404), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[30] ), 
	.D(n6405), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[29] ), 
	.D(n6406), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[28] ), 
	.D(n6407), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[27] ), 
	.D(n6408), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[26] ), 
	.D(n6409), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[25] ), 
	.D(n6410), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[24] ), 
	.D(n6411), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[23] ), 
	.D(n6412), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[22] ), 
	.D(n6413), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[21] ), 
	.D(n6414), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[20] ), 
	.D(n6415), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[19] ), 
	.D(n6416), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[18] ), 
	.D(n6417), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[17] ), 
	.D(n6418), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[16] ), 
	.D(n6419), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[15] ), 
	.D(n6420), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[14] ), 
	.D(n6421), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[13] ), 
	.D(n6422), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[12] ), 
	.D(n6423), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[11] ), 
	.D(n6424), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[10] ), 
	.D(n6425), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[9] ), 
	.D(n6426), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[8] ), 
	.D(n6427), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[7] ), 
	.D(n6428), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[6] ), 
	.D(n6429), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[5] ), 
	.D(n6430), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[4] ), 
	.D(n6431), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[3] ), 
	.D(n6432), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[2] ), 
	.D(n6433), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[1] ), 
	.D(n6434), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell10/sr_out[0] ), 
	.D(n6435), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[31] ), 
	.D(n6370), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[30] ), 
	.D(n6371), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[29] ), 
	.D(n6372), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[28] ), 
	.D(n6373), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[27] ), 
	.D(n6374), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[26] ), 
	.D(n6375), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[25] ), 
	.D(n6376), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[24] ), 
	.D(n6377), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[23] ), 
	.D(n6378), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[22] ), 
	.D(n6379), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[21] ), 
	.D(n6380), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[20] ), 
	.D(n6381), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[19] ), 
	.D(n6382), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[18] ), 
	.D(n6383), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[17] ), 
	.D(n6384), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[16] ), 
	.D(n6385), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[15] ), 
	.D(n6386), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[14] ), 
	.D(n6387), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[13] ), 
	.D(n6388), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[12] ), 
	.D(n6389), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[11] ), 
	.D(n6390), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[10] ), 
	.D(n6391), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[9] ), 
	.D(n6392), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[8] ), 
	.D(n6393), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[7] ), 
	.D(n6394), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[6] ), 
	.D(n6395), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[5] ), 
	.D(n6396), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[4] ), 
	.D(n6397), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[3] ), 
	.D(n6398), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[2] ), 
	.D(n6399), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[1] ), 
	.D(n6400), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell11/sr_out[0] ), 
	.D(n6401), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[31] ), 
	.D(n6336), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[30] ), 
	.D(n6337), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[29] ), 
	.D(n6338), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[28] ), 
	.D(n6339), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[27] ), 
	.D(n6340), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[26] ), 
	.D(n6341), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[25] ), 
	.D(n6342), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[24] ), 
	.D(n6343), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[23] ), 
	.D(n6344), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[22] ), 
	.D(n6345), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[21] ), 
	.D(n6346), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[20] ), 
	.D(n6347), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[19] ), 
	.D(n6348), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[18] ), 
	.D(n6349), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[17] ), 
	.D(n6350), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[16] ), 
	.D(n6351), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[15] ), 
	.D(n6352), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[14] ), 
	.D(n6353), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[13] ), 
	.D(n6354), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[12] ), 
	.D(n6355), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[11] ), 
	.D(n6356), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[10] ), 
	.D(n6357), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[9] ), 
	.D(n6358), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[8] ), 
	.D(n6359), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[7] ), 
	.D(n6360), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[6] ), 
	.D(n6361), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[5] ), 
	.D(n6362), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[4] ), 
	.D(n6363), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[3] ), 
	.D(n6364), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[2] ), 
	.D(n6365), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[1] ), 
	.D(n6366), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell12/sr_out[0] ), 
	.D(n6367), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[31] ), 
	.D(n6302), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[30] ), 
	.D(n6303), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[29] ), 
	.D(n6304), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[28] ), 
	.D(n6305), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[27] ), 
	.D(n6306), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[26] ), 
	.D(n6307), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[25] ), 
	.D(n6308), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[24] ), 
	.D(n6309), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[23] ), 
	.D(n6310), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[22] ), 
	.D(n6311), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[21] ), 
	.D(n6312), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[20] ), 
	.D(n6313), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[19] ), 
	.D(n6314), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[18] ), 
	.D(n6315), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[17] ), 
	.D(n6316), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[16] ), 
	.D(n6317), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[15] ), 
	.D(n6318), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[14] ), 
	.D(n6319), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[13] ), 
	.D(n6320), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[12] ), 
	.D(n6321), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[11] ), 
	.D(n6322), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[10] ), 
	.D(n6323), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[9] ), 
	.D(n6324), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[8] ), 
	.D(n6325), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[7] ), 
	.D(n6326), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[6] ), 
	.D(n6327), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[5] ), 
	.D(n6328), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[4] ), 
	.D(n6329), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[3] ), 
	.D(n6330), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[2] ), 
	.D(n6331), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[1] ), 
	.D(n6332), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell13/sr_out[0] ), 
	.D(n6333), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[31] ), 
	.D(n6268), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[30] ), 
	.D(n6269), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[29] ), 
	.D(n6270), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[28] ), 
	.D(n6271), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[27] ), 
	.D(n6272), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[26] ), 
	.D(n6273), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[25] ), 
	.D(n6274), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[24] ), 
	.D(n6275), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[23] ), 
	.D(n6276), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[22] ), 
	.D(n6277), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[21] ), 
	.D(n6278), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[20] ), 
	.D(n6279), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[19] ), 
	.D(n6280), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[18] ), 
	.D(n6281), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[17] ), 
	.D(n6282), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[16] ), 
	.D(n6283), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[15] ), 
	.D(n6284), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[14] ), 
	.D(n6285), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[13] ), 
	.D(n6286), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[12] ), 
	.D(n6287), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[11] ), 
	.D(n6288), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[10] ), 
	.D(n6289), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[9] ), 
	.D(n6290), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[8] ), 
	.D(n6291), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[7] ), 
	.D(n6292), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[6] ), 
	.D(n6293), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[5] ), 
	.D(n6294), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[4] ), 
	.D(n6295), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[3] ), 
	.D(n6296), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[2] ), 
	.D(n6297), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[1] ), 
	.D(n6298), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell14/sr_out[0] ), 
	.D(n6299), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[31]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[31] ), 
	.D(n6234), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[30]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[30] ), 
	.D(n6235), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[29]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[29] ), 
	.D(n6236), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[28]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[28] ), 
	.D(n6237), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[27]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[27] ), 
	.D(n6238), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[26]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[26] ), 
	.D(n6239), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[25]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[25] ), 
	.D(n6240), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[24]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[24] ), 
	.D(n6241), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[23]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[23] ), 
	.D(n6242), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[22]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[22] ), 
	.D(n6243), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[21]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[21] ), 
	.D(n6244), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[20]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[20] ), 
	.D(n6245), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[19]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[19] ), 
	.D(n6246), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[18]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[18] ), 
	.D(n6247), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[17]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[17] ), 
	.D(n6248), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[16]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[16] ), 
	.D(n6249), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[15]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[15] ), 
	.D(n6250), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[14]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[14] ), 
	.D(n6251), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[13]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[13] ), 
	.D(n6252), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[12]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[12] ), 
	.D(n6253), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[11]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[11] ), 
	.D(n6254), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[10]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[10] ), 
	.D(n6255), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[9]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[9] ), 
	.D(n6256), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[8]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[8] ), 
	.D(n6257), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[7]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[7] ), 
	.D(n6258), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[6]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[6] ), 
	.D(n6259), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[5]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[5] ), 
	.D(n6260), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[4]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[4] ), 
	.D(n6261), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[3]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[3] ), 
	.D(n6262), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[2]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[2] ), 
	.D(n6263), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[1]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[1] ), 
	.D(n6264), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/register/sr_reg[0]  (.Q(\fifo_from_fir/fifo_cell15/sr_out[0] ), 
	.D(n6265), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[31] ), 
	.D(n5420), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[30] ), 
	.D(n5421), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[29] ), 
	.D(n5422), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[28] ), 
	.D(n5423), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[27] ), 
	.D(n5424), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[26] ), 
	.D(n5425), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[25] ), 
	.D(n5426), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[24] ), 
	.D(n5427), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[23] ), 
	.D(n5428), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[22] ), 
	.D(n5429), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[21] ), 
	.D(n5430), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[20] ), 
	.D(n5431), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[19] ), 
	.D(n5432), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[18] ), 
	.D(n5433), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[17] ), 
	.D(n5434), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[16] ), 
	.D(n5435), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[15] ), 
	.D(n5436), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[14] ), 
	.D(n5437), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[13] ), 
	.D(n5438), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[12] ), 
	.D(n5439), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[11] ), 
	.D(n5440), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[10] ), 
	.D(n5441), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[9] ), 
	.D(n5442), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[8] ), 
	.D(n5443), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[7] ), 
	.D(n5444), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[6] ), 
	.D(n5445), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[5] ), 
	.D(n5446), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[4] ), 
	.D(n5447), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[3] ), 
	.D(n5448), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[2] ), 
	.D(n5449), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[1] ), 
	.D(n5450), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell0/sr_out[0] ), 
	.D(n5451), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[31] ), 
	.D(n6181), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[30] ), 
	.D(n6182), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[29] ), 
	.D(n6183), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[28] ), 
	.D(n6184), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[27] ), 
	.D(n6185), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[26] ), 
	.D(n6186), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[25] ), 
	.D(n6187), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[24] ), 
	.D(n6188), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[23] ), 
	.D(n6189), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[22] ), 
	.D(n6190), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[21] ), 
	.D(n6191), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[20] ), 
	.D(n6192), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[19] ), 
	.D(n6193), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[18] ), 
	.D(n6194), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[17] ), 
	.D(n6195), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[16] ), 
	.D(n6196), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[15] ), 
	.D(n6197), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[14] ), 
	.D(n6198), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[13] ), 
	.D(n6199), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[12] ), 
	.D(n6200), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[11] ), 
	.D(n6201), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[10] ), 
	.D(n6202), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[9] ), 
	.D(n6203), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[8] ), 
	.D(n6204), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[7] ), 
	.D(n6205), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[6] ), 
	.D(n6206), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[5] ), 
	.D(n6207), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[4] ), 
	.D(n6208), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[3] ), 
	.D(n6209), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[2] ), 
	.D(n6210), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[1] ), 
	.D(n6211), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell1/sr_out[0] ), 
	.D(n6212), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[31] ), 
	.D(n6147), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[30] ), 
	.D(n6148), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[29] ), 
	.D(n6149), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[28] ), 
	.D(n6150), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[27] ), 
	.D(n6151), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[26] ), 
	.D(n6152), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[25] ), 
	.D(n6153), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[24] ), 
	.D(n6154), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[23] ), 
	.D(n6155), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[22] ), 
	.D(n6156), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[21] ), 
	.D(n6157), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[20] ), 
	.D(n6158), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[19] ), 
	.D(n6159), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[18] ), 
	.D(n6160), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[17] ), 
	.D(n6161), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[16] ), 
	.D(n6162), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[15] ), 
	.D(n6163), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[14] ), 
	.D(n6164), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[13] ), 
	.D(n6165), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[12] ), 
	.D(n6166), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[11] ), 
	.D(n6167), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[10] ), 
	.D(n6168), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[9] ), 
	.D(n6169), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[8] ), 
	.D(n6170), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[7] ), 
	.D(n6171), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[6] ), 
	.D(n6172), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[5] ), 
	.D(n6173), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[4] ), 
	.D(n6174), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[3] ), 
	.D(n6175), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[2] ), 
	.D(n6176), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[1] ), 
	.D(n6177), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell2/sr_out[0] ), 
	.D(n6178), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[31] ), 
	.D(n6113), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[30] ), 
	.D(n6114), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[29] ), 
	.D(n6115), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[28] ), 
	.D(n6116), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[27] ), 
	.D(n6117), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[26] ), 
	.D(n6118), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[25] ), 
	.D(n6119), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[24] ), 
	.D(n6120), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[23] ), 
	.D(n6121), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[22] ), 
	.D(n6122), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[21] ), 
	.D(n6123), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[20] ), 
	.D(n6124), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[19] ), 
	.D(n6125), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[18] ), 
	.D(n6126), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[17] ), 
	.D(n6127), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[16] ), 
	.D(n6128), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[15] ), 
	.D(n6129), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[14] ), 
	.D(n6130), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[13] ), 
	.D(n6131), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[12] ), 
	.D(n6132), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[11] ), 
	.D(n6133), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[10] ), 
	.D(n6134), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[9] ), 
	.D(n6135), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[8] ), 
	.D(n6136), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[7] ), 
	.D(n6137), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[6] ), 
	.D(n6138), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[5] ), 
	.D(n6139), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[4] ), 
	.D(n6140), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[3] ), 
	.D(n6141), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[2] ), 
	.D(n6142), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[1] ), 
	.D(n6143), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell3/sr_out[0] ), 
	.D(n6144), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[31] ), 
	.D(n6079), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[30] ), 
	.D(n6080), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[29] ), 
	.D(n6081), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[28] ), 
	.D(n6082), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[27] ), 
	.D(n6083), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[26] ), 
	.D(n6084), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[25] ), 
	.D(n6085), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[24] ), 
	.D(n6086), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[23] ), 
	.D(n6087), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[22] ), 
	.D(n6088), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[21] ), 
	.D(n6089), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[20] ), 
	.D(n6090), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[19] ), 
	.D(n6091), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[18] ), 
	.D(n6092), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[17] ), 
	.D(n6093), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[16] ), 
	.D(n6094), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[15] ), 
	.D(n6095), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[14] ), 
	.D(n6096), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[13] ), 
	.D(n6097), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[12] ), 
	.D(n6098), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[11] ), 
	.D(n6099), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[10] ), 
	.D(n6100), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[9] ), 
	.D(n6101), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[8] ), 
	.D(n6102), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[7] ), 
	.D(n6103), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[6] ), 
	.D(n6104), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[5] ), 
	.D(n6105), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[4] ), 
	.D(n6106), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[3] ), 
	.D(n6107), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[2] ), 
	.D(n6108), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[1] ), 
	.D(n6109), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell4/sr_out[0] ), 
	.D(n6110), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[31] ), 
	.D(n6045), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[30] ), 
	.D(n6046), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[29] ), 
	.D(n6047), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[28] ), 
	.D(n6048), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[27] ), 
	.D(n6049), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[26] ), 
	.D(n6050), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[25] ), 
	.D(n6051), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[24] ), 
	.D(n6052), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[23] ), 
	.D(n6053), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[22] ), 
	.D(n6054), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[21] ), 
	.D(n6055), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[20] ), 
	.D(n6056), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[19] ), 
	.D(n6057), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[18] ), 
	.D(n6058), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[17] ), 
	.D(n6059), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[16] ), 
	.D(n6060), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[15] ), 
	.D(n6061), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[14] ), 
	.D(n6062), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[13] ), 
	.D(n6063), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[12] ), 
	.D(n6064), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[11] ), 
	.D(n6065), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[10] ), 
	.D(n6066), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[9] ), 
	.D(n6067), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[8] ), 
	.D(n6068), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[7] ), 
	.D(n6069), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[6] ), 
	.D(n6070), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[5] ), 
	.D(n6071), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[4] ), 
	.D(n6072), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[3] ), 
	.D(n6073), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[2] ), 
	.D(n6074), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[1] ), 
	.D(n6075), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell5/sr_out[0] ), 
	.D(n6076), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[31] ), 
	.D(n6011), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[30] ), 
	.D(n6012), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[29] ), 
	.D(n6013), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[28] ), 
	.D(n6014), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[27] ), 
	.D(n6015), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[26] ), 
	.D(n6016), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[25] ), 
	.D(n6017), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[24] ), 
	.D(n6018), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[23] ), 
	.D(n6019), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[22] ), 
	.D(n6020), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[21] ), 
	.D(n6021), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[20] ), 
	.D(n6022), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[19] ), 
	.D(n6023), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[18] ), 
	.D(n6024), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[17] ), 
	.D(n6025), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[16] ), 
	.D(n6026), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[15] ), 
	.D(n6027), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[14] ), 
	.D(n6028), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[13] ), 
	.D(n6029), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[12] ), 
	.D(n6030), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[11] ), 
	.D(n6031), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[10] ), 
	.D(n6032), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[9] ), 
	.D(n6033), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[8] ), 
	.D(n6034), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[7] ), 
	.D(n6035), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[6] ), 
	.D(n6036), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[5] ), 
	.D(n6037), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[4] ), 
	.D(n6038), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[3] ), 
	.D(n6039), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[2] ), 
	.D(n6040), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[1] ), 
	.D(n6041), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell6/sr_out[0] ), 
	.D(n6042), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[31] ), 
	.D(n5977), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[30] ), 
	.D(n5978), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[29] ), 
	.D(n5979), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[28] ), 
	.D(n5980), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[27] ), 
	.D(n5981), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[26] ), 
	.D(n5982), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[25] ), 
	.D(n5983), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[24] ), 
	.D(n5984), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[23] ), 
	.D(n5985), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[22] ), 
	.D(n5986), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[21] ), 
	.D(n5987), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[20] ), 
	.D(n5988), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[19] ), 
	.D(n5989), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[18] ), 
	.D(n5990), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[17] ), 
	.D(n5991), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[16] ), 
	.D(n5992), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[15] ), 
	.D(n5993), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[14] ), 
	.D(n5994), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[13] ), 
	.D(n5995), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[12] ), 
	.D(n5996), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[11] ), 
	.D(n5997), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[10] ), 
	.D(n5998), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[9] ), 
	.D(n5999), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[8] ), 
	.D(n6000), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[7] ), 
	.D(n6001), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[6] ), 
	.D(n6002), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[5] ), 
	.D(n6003), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[4] ), 
	.D(n6004), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[3] ), 
	.D(n6005), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[2] ), 
	.D(n6006), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[1] ), 
	.D(n6007), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell7/sr_out[0] ), 
	.D(n6008), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[31] ), 
	.D(n5943), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[30] ), 
	.D(n5944), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[29] ), 
	.D(n5945), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[28] ), 
	.D(n5946), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[27] ), 
	.D(n5947), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[26] ), 
	.D(n5948), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[25] ), 
	.D(n5949), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[24] ), 
	.D(n5950), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[23] ), 
	.D(n5951), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[22] ), 
	.D(n5952), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[21] ), 
	.D(n5953), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[20] ), 
	.D(n5954), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[19] ), 
	.D(n5955), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[18] ), 
	.D(n5956), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[17] ), 
	.D(n5957), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[16] ), 
	.D(n5958), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[15] ), 
	.D(n5959), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[14] ), 
	.D(n5960), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[13] ), 
	.D(n5961), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[12] ), 
	.D(n5962), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[11] ), 
	.D(n5963), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[10] ), 
	.D(n5964), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[9] ), 
	.D(n5965), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[8] ), 
	.D(n5966), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[7] ), 
	.D(n5967), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[6] ), 
	.D(n5968), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[5] ), 
	.D(n5969), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[4] ), 
	.D(n5970), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[3] ), 
	.D(n5971), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[2] ), 
	.D(n5972), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[1] ), 
	.D(n5973), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell8/sr_out[0] ), 
	.D(n5974), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[31] ), 
	.D(n5909), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[30] ), 
	.D(n5910), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[29] ), 
	.D(n5911), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[28] ), 
	.D(n5912), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[27] ), 
	.D(n5913), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[26] ), 
	.D(n5914), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[25] ), 
	.D(n5915), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[24] ), 
	.D(n5916), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[23] ), 
	.D(n5917), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[22] ), 
	.D(n5918), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[21] ), 
	.D(n5919), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[20] ), 
	.D(n5920), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[19] ), 
	.D(n5921), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[18] ), 
	.D(n5922), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[17] ), 
	.D(n5923), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[16] ), 
	.D(n5924), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[15] ), 
	.D(n5925), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[14] ), 
	.D(n5926), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[13] ), 
	.D(n5927), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[12] ), 
	.D(n5928), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[11] ), 
	.D(n5929), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[10] ), 
	.D(n5930), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[9] ), 
	.D(n5931), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[8] ), 
	.D(n5932), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[7] ), 
	.D(n5933), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[6] ), 
	.D(n5934), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[5] ), 
	.D(n5935), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[4] ), 
	.D(n5936), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[3] ), 
	.D(n5937), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[2] ), 
	.D(n5938), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[1] ), 
	.D(n5939), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell9/sr_out[0] ), 
	.D(n5940), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[31] ), 
	.D(n5875), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[30] ), 
	.D(n5876), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[29] ), 
	.D(n5877), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[28] ), 
	.D(n5878), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[27] ), 
	.D(n5879), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[26] ), 
	.D(n5880), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[25] ), 
	.D(n5881), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[24] ), 
	.D(n5882), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[23] ), 
	.D(n5883), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[22] ), 
	.D(n5884), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[21] ), 
	.D(n5885), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[20] ), 
	.D(n5886), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[19] ), 
	.D(n5887), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[18] ), 
	.D(n5888), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[17] ), 
	.D(n5889), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[16] ), 
	.D(n5890), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[15] ), 
	.D(n5891), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[14] ), 
	.D(n5892), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[13] ), 
	.D(n5893), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[12] ), 
	.D(n5894), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[11] ), 
	.D(n5895), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[10] ), 
	.D(n5896), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[9] ), 
	.D(n5897), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[8] ), 
	.D(n5898), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[7] ), 
	.D(n5899), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[6] ), 
	.D(n5900), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[5] ), 
	.D(n5901), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[4] ), 
	.D(n5902), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[3] ), 
	.D(n5903), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[2] ), 
	.D(n5904), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[1] ), 
	.D(n5905), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell10/sr_out[0] ), 
	.D(n5906), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[31] ), 
	.D(n5841), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[30] ), 
	.D(n5842), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[29] ), 
	.D(n5843), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[28] ), 
	.D(n5844), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[27] ), 
	.D(n5845), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[26] ), 
	.D(n5846), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[25] ), 
	.D(n5847), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[24] ), 
	.D(n5848), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[23] ), 
	.D(n5849), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[22] ), 
	.D(n5850), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[21] ), 
	.D(n5851), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[20] ), 
	.D(n5852), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[19] ), 
	.D(n5853), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[18] ), 
	.D(n5854), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[17] ), 
	.D(n5855), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[16] ), 
	.D(n5856), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[15] ), 
	.D(n5857), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[14] ), 
	.D(n5858), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[13] ), 
	.D(n5859), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[12] ), 
	.D(n5860), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[11] ), 
	.D(n5861), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[10] ), 
	.D(n5862), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[9] ), 
	.D(n5863), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[8] ), 
	.D(n5864), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[7] ), 
	.D(n5865), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[6] ), 
	.D(n5866), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[5] ), 
	.D(n5867), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[4] ), 
	.D(n5868), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[3] ), 
	.D(n5869), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[2] ), 
	.D(n5870), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[1] ), 
	.D(n5871), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell11/sr_out[0] ), 
	.D(n5872), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[31] ), 
	.D(n5807), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[30] ), 
	.D(n5808), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[29] ), 
	.D(n5809), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[28] ), 
	.D(n5810), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[27] ), 
	.D(n5811), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[26] ), 
	.D(n5812), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[25] ), 
	.D(n5813), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[24] ), 
	.D(n5814), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[23] ), 
	.D(n5815), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[22] ), 
	.D(n5816), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[21] ), 
	.D(n5817), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[20] ), 
	.D(n5818), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[19] ), 
	.D(n5819), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[18] ), 
	.D(n5820), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[17] ), 
	.D(n5821), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[16] ), 
	.D(n5822), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[15] ), 
	.D(n5823), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[14] ), 
	.D(n5824), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[13] ), 
	.D(n5825), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[12] ), 
	.D(n5826), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[11] ), 
	.D(n5827), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[10] ), 
	.D(n5828), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[9] ), 
	.D(n5829), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[8] ), 
	.D(n5830), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[7] ), 
	.D(n5831), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[6] ), 
	.D(n5832), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[5] ), 
	.D(n5833), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[4] ), 
	.D(n5834), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[3] ), 
	.D(n5835), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[2] ), 
	.D(n5836), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[1] ), 
	.D(n5837), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell12/sr_out[0] ), 
	.D(n5838), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[31] ), 
	.D(n5773), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[30] ), 
	.D(n5774), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[29] ), 
	.D(n5775), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[28] ), 
	.D(n5776), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[27] ), 
	.D(n5777), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[26] ), 
	.D(n5778), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[25] ), 
	.D(n5779), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[24] ), 
	.D(n5780), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[23] ), 
	.D(n5781), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[22] ), 
	.D(n5782), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[21] ), 
	.D(n5783), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[20] ), 
	.D(n5784), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[19] ), 
	.D(n5785), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[18] ), 
	.D(n5786), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[17] ), 
	.D(n5787), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[16] ), 
	.D(n5788), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[15] ), 
	.D(n5789), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[14] ), 
	.D(n5790), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[13] ), 
	.D(n5791), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[12] ), 
	.D(n5792), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[11] ), 
	.D(n5793), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[10] ), 
	.D(n5794), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[9] ), 
	.D(n5795), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[8] ), 
	.D(n5796), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[7] ), 
	.D(n5797), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[6] ), 
	.D(n5798), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[5] ), 
	.D(n5799), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[4] ), 
	.D(n5800), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[3] ), 
	.D(n5801), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[2] ), 
	.D(n5802), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[1] ), 
	.D(n5803), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell13/sr_out[0] ), 
	.D(n5804), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[31] ), 
	.D(n5739), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[30] ), 
	.D(n5740), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[29] ), 
	.D(n5741), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[28] ), 
	.D(n5742), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[27] ), 
	.D(n5743), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[26] ), 
	.D(n5744), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[25] ), 
	.D(n5745), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[24] ), 
	.D(n5746), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[23] ), 
	.D(n5747), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[22] ), 
	.D(n5748), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[21] ), 
	.D(n5749), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[20] ), 
	.D(n5750), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[19] ), 
	.D(n5751), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[18] ), 
	.D(n5752), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[17] ), 
	.D(n5753), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[16] ), 
	.D(n5754), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[15] ), 
	.D(n5755), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[14] ), 
	.D(n5756), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[13] ), 
	.D(n5757), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[12] ), 
	.D(n5758), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[11] ), 
	.D(n5759), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[10] ), 
	.D(n5760), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[9] ), 
	.D(n5761), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[8] ), 
	.D(n5762), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[7] ), 
	.D(n5763), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[6] ), 
	.D(n5764), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[5] ), 
	.D(n5765), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[4] ), 
	.D(n5766), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[3] ), 
	.D(n5767), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[2] ), 
	.D(n5768), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[1] ), 
	.D(n5769), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell14/sr_out[0] ), 
	.D(n5770), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[31]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[31] ), 
	.D(n5705), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[30]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[30] ), 
	.D(n5706), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[29]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[29] ), 
	.D(n5707), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[28]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[28] ), 
	.D(n5708), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[27]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[27] ), 
	.D(n5709), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[26]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[26] ), 
	.D(n5710), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[25]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[25] ), 
	.D(n5711), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[24]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[24] ), 
	.D(n5712), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[23]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[23] ), 
	.D(n5713), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[22]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[22] ), 
	.D(n5714), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[21]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[21] ), 
	.D(n5715), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[20]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[20] ), 
	.D(n5716), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[19]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[19] ), 
	.D(n5717), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[18]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[18] ), 
	.D(n5718), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[17]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[17] ), 
	.D(n5719), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[16]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[16] ), 
	.D(n5720), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[15]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[15] ), 
	.D(n5721), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[14]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[14] ), 
	.D(n5722), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[13]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[13] ), 
	.D(n5723), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[12]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[12] ), 
	.D(n5724), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[11]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[11] ), 
	.D(n5725), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[10]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[10] ), 
	.D(n5726), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[9]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[9] ), 
	.D(n5727), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[8]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[8] ), 
	.D(n5728), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[7]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[7] ), 
	.D(n5729), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[6]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[6] ), 
	.D(n5730), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[5]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[5] ), 
	.D(n5731), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[4]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[4] ), 
	.D(n5732), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[3]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[3] ), 
	.D(n5733), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[2]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[2] ), 
	.D(n5734), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[1]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[1] ), 
	.D(n5735), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/register/sr_reg[0]  (.Q(\fifo_from_fft/fifo_cell15/sr_out[0] ), 
	.D(n5736), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fir/fifo_cell0/controller/write_enable_reg  (.RN(n9546), 
	.QN(\fifo_from_fir/fifo_cell0/controller/write_enable ), 
	.E(\fifo_from_fir/fifo_cell0/controller/valid_read ), 
	.D(n7216), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \fifo_from_fft/fifo_cell0/controller/write_enable_reg  (.RN(n9546), 
	.QN(\fifo_from_fft/fifo_cell0/controller/write_enable ), 
	.E(\fifo_from_fft/fifo_cell0/controller/valid_read ), 
	.D(n7221), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/pla_top/instruction_valid_reg  (.Q(\router/pla_top/instruction_valid ), 
	.D(\router/pla_top/N60 ), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell15/reg_gtok/token ), 
	.D(n6745), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell15/reg_gtok/token ), 
	.D(n6216), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell15/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell15/reg_gtok/token ), 
	.D(n5469), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell15/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell15/reg_gtok/token ), 
	.D(n5521), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell0/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell0/controller/valid_read ), 
	.D(n9515), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell0/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell0/controller/valid_read ), 
	.D(n9524), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell0/controller/valid_read ), 
	.D(n9520), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell0/controller/valid_read ), 
	.D(n9528), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell15/reg_ptok/token_reg  (.Q(\fifo_to_fft/hang[14] ), 
	.D(n5516), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell15/reg_ptok/token_reg  (.Q(\fifo_to_fir/hang[14] ), 
	.D(n5568), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/iir_write_calc/counter/hold_reg  (.Q(\router/addr_calc/iir_write_calc/counter/hold ), 
	.D(n6766), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/fir_read_calc/counter/hold_reg  (.Q(\router/addr_calc/fir_read_calc/counter/hold ), 
	.D(n5572), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/fir_write_calc/counter/hold_reg  (.Q(\router/addr_calc/fir_write_calc/counter/hold ), 
	.D(n5520), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/fft_read_calc/counter/hold_reg  (.Q(\router/addr_calc/fft_read_calc/counter/hold ), 
	.D(n5457), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/fft_write_calc/counter/hold_reg  (.Q(\router/addr_calc/fft_write_calc/counter/hold ), 
	.D(n5468), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/data_out/en_reg  (.Q(\fifo_from_fir/fifo_cell0/data_out/N9 ), 
	.D(n4766), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/data_out/en_reg  (.Q(\fifo_from_fft/fifo_cell0/data_out/N9 ), 
	.D(n4580), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell14/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell13/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell14/data_out/N9 ), 
	.Q(n8093), 
	.D(FE_OFN735_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell13/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell12/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell13/data_out/N9 ), 
	.Q(n8092), 
	.D(FE_OFN736_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell12/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell11/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell12/data_out/N9 ), 
	.Q(n8091), 
	.D(FE_OFN736_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell11/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell10/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell11/data_out/N9 ), 
	.Q(n8090), 
	.D(FE_OFN739_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell10/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell9/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell10/data_out/N9 ), 
	.Q(n8089), 
	.D(FE_OFN737_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell9/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell8/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell9/data_out/N9 ), 
	.Q(n8088), 
	.D(FE_OFN744_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell8/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell7/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell8/data_out/N9 ), 
	.Q(n8087), 
	.D(FE_OFN744_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell7/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell6/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell7/data_out/N9 ), 
	.Q(n8086), 
	.D(FE_OFN743_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell6/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell5/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell6/data_out/N9 ), 
	.Q(n8085), 
	.D(FE_OFN740_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell5/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell4/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell5/data_out/N9 ), 
	.Q(n8084), 
	.D(FE_OFN740_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell4/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell3/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell4/data_out/N9 ), 
	.Q(n8083), 
	.D(FE_OFN738_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell3/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell2/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell3/data_out/N9 ), 
	.Q(n8082), 
	.D(FE_OFN736_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell2/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell1/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell2/data_out/N9 ), 
	.Q(n8081), 
	.D(n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell1/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell0/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell1/data_out/N9 ), 
	.Q(n8080), 
	.D(FE_OFN735_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell14/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell13/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell14/data_out/N9 ), 
	.Q(n8078), 
	.D(FE_OFN723_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell13/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell12/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell13/data_out/N9 ), 
	.Q(n8077), 
	.D(FE_OFN722_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell12/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell11/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell12/data_out/N9 ), 
	.Q(n8076), 
	.D(FE_OFN728_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell11/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell10/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell11/data_out/N9 ), 
	.Q(n8075), 
	.D(FE_OFN725_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell10/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell9/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell10/data_out/N9 ), 
	.Q(n8074), 
	.D(FE_OFN726_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell9/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell8/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell9/data_out/N9 ), 
	.Q(n8073), 
	.D(FE_OFN728_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell8/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell7/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell8/data_out/N9 ), 
	.Q(n8072), 
	.D(FE_OFN727_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell7/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell6/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell7/data_out/N9 ), 
	.Q(n8071), 
	.D(FE_OFN722_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell6/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell5/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell6/data_out/N9 ), 
	.Q(n8070), 
	.D(FE_OFN1822_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell5/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell4/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell5/data_out/N9 ), 
	.Q(n8069), 
	.D(FE_OFN1822_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell4/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell3/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell4/data_out/N9 ), 
	.Q(n8068), 
	.D(FE_OFN1823_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell3/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell2/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell3/data_out/N9 ), 
	.Q(n8067), 
	.D(FE_OFN1822_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell2/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell1/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell2/data_out/N9 ), 
	.Q(n8066), 
	.D(FE_OFN1822_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell1/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell0/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell1/data_out/N9 ), 
	.Q(n8065), 
	.D(FE_OFN720_n4643), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell15/data_out/en_reg  (.RN(\fifo_from_fir/fifo_cell14/reg_gtok/token ), 
	.QN(\fifo_from_fir/fifo_cell15/data_out/N9 ), 
	.Q(n8094), 
	.D(FE_OFN741_n4829), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell15/data_out/en_reg  (.RN(\fifo_from_fft/fifo_cell14/reg_gtok/token ), 
	.QN(\fifo_from_fft/fifo_cell15/data_out/N9 ), 
	.Q(n8079), 
	.D(FE_OFN724_n4643), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[31]  (.Q(\router/data_cntl/data_in[31] ), 
	.D(n5351), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[30]  (.Q(\router/data_cntl/data_in[30] ), 
	.D(n5352), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[29]  (.Q(\router/data_cntl/data_in[29] ), 
	.D(n5353), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[28]  (.Q(\router/data_cntl/data_in[28] ), 
	.D(n5354), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[27]  (.Q(\router/data_cntl/data_in[27] ), 
	.D(n5355), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[26]  (.Q(\router/data_cntl/data_in[26] ), 
	.D(n5356), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[25]  (.Q(\router/data_cntl/data_in[25] ), 
	.D(n5357), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[24]  (.Q(\router/data_cntl/data_in[24] ), 
	.D(n5358), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[23]  (.Q(\router/data_cntl/data_in[23] ), 
	.D(n5359), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[22]  (.Q(\router/data_cntl/data_in[22] ), 
	.D(n5360), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[21]  (.Q(\router/data_cntl/data_in[21] ), 
	.D(n5361), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[20]  (.Q(\router/data_cntl/data_in[20] ), 
	.D(n5362), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[19]  (.Q(\router/data_cntl/data_in[19] ), 
	.D(n5363), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[18]  (.Q(\router/data_cntl/data_in[18] ), 
	.D(n5364), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[17]  (.Q(\router/data_cntl/data_in[17] ), 
	.D(n5365), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[16]  (.Q(\router/data_cntl/data_in[16] ), 
	.D(n5366), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[15]  (.Q(\router/data_cntl/data_in[15] ), 
	.D(n5367), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[14]  (.Q(\router/data_cntl/data_in[14] ), 
	.D(n5368), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[13]  (.Q(\router/data_cntl/data_in[13] ), 
	.D(n5369), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[12]  (.Q(\router/data_cntl/data_in[12] ), 
	.D(n5370), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[11]  (.Q(\router/data_cntl/data_in[11] ), 
	.D(n5371), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[10]  (.Q(\router/data_cntl/data_in[10] ), 
	.D(n5372), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[9]  (.Q(\router/data_cntl/data_in[9] ), 
	.D(n5373), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[8]  (.Q(\router/data_cntl/data_in[8] ), 
	.D(n5374), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[7]  (.Q(\router/data_cntl/data_in[7] ), 
	.D(n5375), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[6]  (.Q(\router/data_cntl/data_in[6] ), 
	.D(n5376), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[5]  (.Q(\router/data_cntl/data_in[5] ), 
	.D(n5377), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[4]  (.Q(\router/data_cntl/data_in[4] ), 
	.D(n5378), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[3]  (.Q(\router/data_cntl/data_in[3] ), 
	.D(n5379), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[2]  (.Q(\router/data_cntl/data_in[2] ), 
	.D(n5380), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[1]  (.Q(\router/data_cntl/data_in[1] ), 
	.D(n5381), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/data_in_reg[0]  (.Q(\router/data_cntl/data_in[0] ), 
	.D(n5382), 
	.CK(clk__L1_N0));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1313_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1313_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1313_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1313_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1310_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1310_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1310_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1014_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1017_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(FE_OFN1017_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1014_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1014_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1016_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1017_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1015_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1017_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1015_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1016_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1015_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1016_n2569), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1311_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1311_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1312_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1312_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1311_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(FE_OFN1312_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell15/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1312_n8094), 
	.A(\fifo_from_fir/fifo_cell15/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1435_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1433_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1435_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1435_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1433_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1433_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1134_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1133_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(FE_OFN1133_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(FE_OFN1134_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1136_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1134_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1136_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1135_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1135_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1137_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1135_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1137_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1135_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1137_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1137_n2505), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1436_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1434_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1434_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1437_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1437_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1436_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(FE_OFN1437_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell14/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1436_n8093), 
	.A(\fifo_from_fir/fifo_cell14/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1432_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1432_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1432_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1432_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1429_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1430_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1430_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1430_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1129_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(FE_OFN1132_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1132_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1132_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1132_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1130_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1129_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1130_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1129_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1131_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1131_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1131_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1131_n2441), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1429_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1429_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1431_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1431_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(FE_OFN1431_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell13/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1431_n8092), 
	.A(\fifo_from_fir/fifo_cell13/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1428_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1428_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1428_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1428_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1427_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1427_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1427_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1427_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1124_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1128_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(FE_OFN1128_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1125_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1124_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1124_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1126_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1128_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1125_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1128_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1127_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1126_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1127_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1127_n2377), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1425_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1425_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1426_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1426_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(FE_OFN1426_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell12/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1426_n8091), 
	.A(\fifo_from_fir/fifo_cell12/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1424_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1424_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1424_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1424_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1422_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1423_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1423_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1423_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1123_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(FE_OFN1120_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1121_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1120_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1120_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1123_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1123_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1121_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1123_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1121_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1122_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1122_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1122_n2313), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1421_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1420_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1422_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1420_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1421_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1421_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell11/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1421_n8090), 
	.A(\fifo_from_fir/fifo_cell11/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1419_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1417_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1419_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1419_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1419_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1418_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1418_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1418_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1115_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1119_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(FE_OFN1115_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1116_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1115_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1116_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1119_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1119_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1116_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1119_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1118_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1117_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1118_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1118_n2249), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1416_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1417_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1418_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1416_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell10/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1416_n8089), 
	.A(\fifo_from_fir/fifo_cell10/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1415_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1415_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1415_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1415_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1414_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1413_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1414_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1414_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1111_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(FE_OFN1111_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(FE_OFN1111_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1112_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1112_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1112_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1113_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1113_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1114_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1113_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1114_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1113_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1114_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1114_n2185), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1412_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1413_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1413_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1412_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1412_n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell9/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(n8088), 
	.A(\fifo_from_fir/fifo_cell9/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1411_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1411_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1411_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1411_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1409_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1409_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1410_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1410_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1108_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1109_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(FE_OFN1106_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(FE_OFN1108_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1107_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1108_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1107_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1106_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1109_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1110_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1109_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1110_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1109_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1110_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1110_n2121), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1407_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1408_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1408_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1408_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1407_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell8/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1407_n8087), 
	.A(\fifo_from_fir/fifo_cell8/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1406_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1406_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1406_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1406_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1405_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1405_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1405_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1405_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1102_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1105_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1103_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1102_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1102_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1105_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1105_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1103_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1105_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1104_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1104_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1104_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1103_n2057), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1403_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1404_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1404_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1403_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1403_n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell7/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(n8086), 
	.A(\fifo_from_fir/fifo_cell7/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1402_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1402_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1402_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1402_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1401_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1400_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1401_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1401_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1097_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1098_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(FE_OFN1098_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(FE_OFN1097_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1099_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1099_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1099_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1100_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1100_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1099_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1098_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1101_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1101_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1101_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1101_n1993), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1399_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1399_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1400_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1400_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1399_n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell6/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(n8085), 
	.A(\fifo_from_fir/fifo_cell6/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1396_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1397_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1397_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1397_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1398_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1398_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1398_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1398_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1093_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1096_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1094_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1093_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1093_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1096_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1096_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1094_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1096_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1094_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1095_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1095_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1095_n1929), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1395_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1396_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1395_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1395_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1394_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1394_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell5/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1394_n8084), 
	.A(\fifo_from_fir/fifo_cell5/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1393_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1391_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1393_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1393_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1391_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1392_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1392_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1392_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1092_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(FE_OFN1089_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1090_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1089_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1089_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1092_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1092_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1090_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1092_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1090_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1091_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1091_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1091_n1865), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1390_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1393_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1390_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1389_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1390_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(FE_OFN1389_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell4/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1389_n8083), 
	.A(\fifo_from_fir/fifo_cell4/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1388_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1388_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1388_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1388_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1387_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1387_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1385_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1385_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1085_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1088_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1086_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1085_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1085_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1088_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1088_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1086_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1088_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1086_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1087_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1087_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1087_n1801), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1384_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1384_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1385_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1384_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1386_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1386_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(FE_OFN1386_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell3/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1386_n8082), 
	.A(\fifo_from_fir/fifo_cell3/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1382_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1382_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1382_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1382_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1380_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1380_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1380_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1083_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(FE_OFN1083_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(FE_OFN1082_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1082_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1082_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1082_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1081_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1083_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1081_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1083_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1084_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1084_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1084_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1084_n1737), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1381_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1381_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1381_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1383_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1383_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(FE_OFN1383_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell2/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1383_n8081), 
	.A(\fifo_from_fir/fifo_cell2/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1379_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1379_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1379_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1379_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1376_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1378_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(FE_OFN1378_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(FE_OFN1378_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1077_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1079_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(FE_OFN1077_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1080_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1078_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1078_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1079_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1078_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1079_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1080_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1079_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1080_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1080_n1673), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1376_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1376_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1377_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1377_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(FE_OFN1377_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell1/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1377_n8080), 
	.A(\fifo_from_fir/fifo_cell1/sr_out[0] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[31]  (.Y(fir_data_in[31]), 
	.OE(FE_OFN1150_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[31] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[30]  (.Y(fir_data_in[30]), 
	.OE(FE_OFN1150_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[30] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[29]  (.Y(fir_data_in[29]), 
	.OE(FE_OFN1150_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[29] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[28]  (.Y(fir_data_in[28]), 
	.OE(FE_OFN1150_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[28] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[27]  (.Y(fir_data_in[27]), 
	.OE(FE_OFN1148_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[27] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[26]  (.Y(fir_data_in[26]), 
	.OE(FE_OFN1148_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[26] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[25]  (.Y(fir_data_in[25]), 
	.OE(n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[25] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[24]  (.Y(fir_data_in[24]), 
	.OE(n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[24] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[23]  (.Y(fir_data_in[23]), 
	.OE(FE_OFN1153_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[23] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[22]  (.Y(fir_data_in[22]), 
	.OE(FE_OFN1154_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[22] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[21]  (.Y(fir_data_in[21]), 
	.OE(FE_OFN1154_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[21] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[20]  (.Y(fir_data_in[20]), 
	.OE(FE_OFN1154_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[20] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[19]  (.Y(fir_data_in[19]), 
	.OE(FE_OFN1153_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[19] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[18]  (.Y(fir_data_in[18]), 
	.OE(FE_OFN1155_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[18] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[17]  (.Y(fir_data_in[17]), 
	.OE(FE_OFN1155_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[17] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[16]  (.Y(fir_data_in[16]), 
	.OE(FE_OFN1155_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[16] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[15]  (.Y(fir_data_in[15]), 
	.OE(FE_OFN1156_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[15] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[14]  (.Y(fir_data_in[14]), 
	.OE(FE_OFN1156_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[14] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[13]  (.Y(fir_data_in[13]), 
	.OE(FE_OFN1157_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[13] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[12]  (.Y(fir_data_in[12]), 
	.OE(FE_OFN1156_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[12] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[11]  (.Y(fir_data_in[11]), 
	.OE(FE_OFN1157_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[11] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[10]  (.Y(fir_data_in[10]), 
	.OE(FE_OFN1156_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[10] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[9]  (.Y(fir_data_in[9]), 
	.OE(FE_OFN1157_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[9] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[8]  (.Y(fir_data_in[8]), 
	.OE(FE_OFN1157_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[8] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[7]  (.Y(fir_data_in[7]), 
	.OE(FE_OFN1149_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[7] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[6]  (.Y(fir_data_in[6]), 
	.OE(FE_OFN1149_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[6] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[5]  (.Y(fir_data_in[5]), 
	.OE(FE_OFN1148_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[5] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[4]  (.Y(fir_data_in[4]), 
	.OE(FE_OFN1151_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[4] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[3]  (.Y(fir_data_in[3]), 
	.OE(FE_OFN1152_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[3] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[2]  (.Y(fir_data_in[2]), 
	.OE(FE_OFN1151_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[2] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[1]  (.Y(fir_data_in[1]), 
	.OE(FE_OFN1152_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[1] ));
   TBUFX2TS \fifo_from_fir/fifo_cell0/data_out/do_tri[0]  (.Y(fir_data_in[0]), 
	.OE(FE_OFN1151_n1609), 
	.A(\fifo_from_fir/fifo_cell0/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1309_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1309_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1309_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1309_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1307_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1308_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1306_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1306_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1009_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1013_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1013_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1009_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1009_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(FE_OFN1011_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(FE_OFN1011_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1010_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1011_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1010_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1011_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1012_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1013_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1012_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1012_n1545), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1307_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1308_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1306_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1307_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell15/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1308_n8079), 
	.A(\fifo_from_fft/fifo_cell15/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1375_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1375_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1375_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1375_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1373_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1373_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1073_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1076_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1076_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1073_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1073_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1074_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1074_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1075_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1074_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1075_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1076_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1076_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1075_n1481), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1372_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1371_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1373_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(FE_OFN1371_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1374_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1372_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1372_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell14/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1374_n8078), 
	.A(\fifo_from_fft/fifo_cell14/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1368_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1367_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1368_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1368_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1369_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1369_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1370_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1370_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1072_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1072_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1072_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1072_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1069_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1070_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1069_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1070_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1069_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1070_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1071_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1071_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1071_n1417), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1366_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1366_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1366_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1369_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1370_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1370_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell13/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1367_n8077), 
	.A(\fifo_from_fft/fifo_cell13/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1365_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1365_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1365_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1365_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1363_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1364_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1065_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1068_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1068_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1065_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(FE_OFN1065_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1065_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1066_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1066_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1067_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1066_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1068_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1068_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1067_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1067_n1353), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1362_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1362_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1362_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1364_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1363_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1363_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell12/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1364_n8076), 
	.A(\fifo_from_fft/fifo_cell12/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1361_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1361_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1361_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1361_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1358_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1360_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1359_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1359_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1061_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1064_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1064_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1061_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1061_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1062_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1062_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1063_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1062_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1064_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1064_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1063_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1063_n1289), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1357_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1357_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(FE_OFN1357_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1360_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1359_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1358_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell11/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1360_n8075), 
	.A(\fifo_from_fft/fifo_cell11/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1356_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1356_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1356_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1356_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1354_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1355_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1353_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1353_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1058_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1060_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1060_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1057_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(FE_OFN1056_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1057_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(FE_OFN1056_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1058_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1057_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1058_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1056_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1059_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1060_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1059_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1059_n1225), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1353_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1355_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1354_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1354_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell10/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1355_n8074), 
	.A(\fifo_from_fft/fifo_cell10/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1352_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1352_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1352_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1352_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1350_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1351_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1052_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1053_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1053_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1052_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(FE_OFN1055_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1055_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1055_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1054_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1055_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1054_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1052_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1053_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1054_n1161), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1349_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1349_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1349_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(FE_OFN1349_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1351_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1350_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1350_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell9/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1351_n8073), 
	.A(\fifo_from_fft/fifo_cell9/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1346_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1345_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1346_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1346_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1347_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1347_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1348_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1348_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1049_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1050_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1050_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1049_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1049_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1048_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1048_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1051_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1048_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1051_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1050_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1051_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1051_n1097), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1344_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1344_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1344_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1347_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1348_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1348_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell8/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1345_n8072), 
	.A(\fifo_from_fft/fifo_cell8/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1343_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1343_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1343_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1343_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1341_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1342_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1339_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1339_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1045_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1047_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1047_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1045_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1045_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(FE_OFN1043_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(FE_OFN1043_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1044_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1044_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1046_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1043_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1046_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1047_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1047_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1046_n1033), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1339_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1341_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1341_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1342_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1340_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1340_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell7/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1342_n8071), 
	.A(\fifo_from_fft/fifo_cell7/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1338_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1338_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1338_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1338_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1336_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1337_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1335_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1335_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1042_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1042_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1042_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1042_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(FE_OFN1039_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1040_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1039_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1040_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1039_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1040_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1041_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1041_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1041_n969), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1335_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1337_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1336_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1336_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell6/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1337_n8070), 
	.A(\fifo_from_fft/fifo_cell6/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1331_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1332_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1332_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1331_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1333_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1333_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1334_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1334_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1035_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1038_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1038_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1035_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(FE_OFN1037_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(FE_OFN1037_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1034_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1037_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1036_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1037_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1036_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1038_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1038_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1036_n905), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1331_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1333_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1334_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1334_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell5/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1332_n8069), 
	.A(\fifo_from_fft/fifo_cell5/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1330_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1330_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1330_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1330_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1328_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1329_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1327_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1030_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1030_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1031_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(FE_OFN1033_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(FE_OFN1033_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1032_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1033_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1032_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1033_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1031_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1030_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1031_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1032_n841), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1328_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1328_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1329_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1327_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1327_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell4/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1329_n8068), 
	.A(\fifo_from_fft/fifo_cell4/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1325_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1326_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1325_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1325_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1324_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1326_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1323_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1323_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1027_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1029_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1029_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1029_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1027_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1026_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1026_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1028_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1026_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1028_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1029_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1028_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1028_n777), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1325_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1326_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1323_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1324_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell3/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1326_n8067), 
	.A(\fifo_from_fft/fifo_cell3/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1319_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1320_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1319_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1319_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1321_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1321_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1322_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1322_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1025_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1025_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1025_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1025_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1022_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1023_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1022_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1023_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1022_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1023_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1024_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1024_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1024_n713), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1318_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1318_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1318_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1320_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1322_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1322_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell2/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1320_n8066), 
	.A(\fifo_from_fft/fifo_cell2/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1317_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1317_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1317_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1317_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1315_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1316_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1314_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1314_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1019_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1021_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1021_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1019_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(FE_OFN1018_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1019_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1018_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1020_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1018_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1020_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1021_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1021_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1020_n649), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1315_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1316_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1314_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1315_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell1/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1316_n8065), 
	.A(\fifo_from_fft/fifo_cell1/sr_out[0] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[31]  (.Y(fft_data_in[31]), 
	.OE(FE_OFN1146_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[31] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[30]  (.Y(fft_data_in[30]), 
	.OE(FE_OFN1145_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[30] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[29]  (.Y(fft_data_in[29]), 
	.OE(FE_OFN1145_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[29] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[28]  (.Y(fft_data_in[28]), 
	.OE(FE_OFN1145_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[28] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[27]  (.Y(fft_data_in[27]), 
	.OE(FE_OFN1140_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[27] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[26]  (.Y(fft_data_in[26]), 
	.OE(FE_OFN1142_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[26] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[25]  (.Y(fft_data_in[25]), 
	.OE(FE_OFN1144_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[25] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[24]  (.Y(fft_data_in[24]), 
	.OE(FE_OFN1144_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[24] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[23]  (.Y(fft_data_in[23]), 
	.OE(FE_OFN1139_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[23] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[22]  (.Y(fft_data_in[22]), 
	.OE(FE_OFN1146_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[22] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[21]  (.Y(fft_data_in[21]), 
	.OE(FE_OFN1146_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[21] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[20]  (.Y(fft_data_in[20]), 
	.OE(FE_OFN1143_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[20] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[19]  (.Y(fft_data_in[19]), 
	.OE(FE_OFN1138_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[19] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[18]  (.Y(fft_data_in[18]), 
	.OE(FE_OFN1138_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[18] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[17]  (.Y(fft_data_in[17]), 
	.OE(FE_OFN1141_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[17] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[16]  (.Y(fft_data_in[16]), 
	.OE(FE_OFN1141_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[16] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[15]  (.Y(fft_data_in[15]), 
	.OE(FE_OFN1143_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[15] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[14]  (.Y(fft_data_in[14]), 
	.OE(FE_OFN1143_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[14] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[13]  (.Y(fft_data_in[13]), 
	.OE(FE_OFN1143_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[13] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[12]  (.Y(fft_data_in[12]), 
	.OE(FE_OFN1141_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[12] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[11]  (.Y(fft_data_in[11]), 
	.OE(FE_OFN1147_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[11] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[10]  (.Y(fft_data_in[10]), 
	.OE(FE_OFN1147_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[10] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[9]  (.Y(fft_data_in[9]), 
	.OE(FE_OFN1147_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[9] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[8]  (.Y(fft_data_in[8]), 
	.OE(FE_OFN1147_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[8] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[7]  (.Y(fft_data_in[7]), 
	.OE(FE_OFN1144_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[7] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[6]  (.Y(fft_data_in[6]), 
	.OE(FE_OFN1139_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[6] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[5]  (.Y(fft_data_in[5]), 
	.OE(FE_OFN1139_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[5] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[4]  (.Y(fft_data_in[4]), 
	.OE(n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[4] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[3]  (.Y(fft_data_in[3]), 
	.OE(FE_OFN1142_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[3] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[2]  (.Y(fft_data_in[2]), 
	.OE(FE_OFN1144_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[2] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[1]  (.Y(fft_data_in[1]), 
	.OE(FE_OFN1140_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[1] ));
   TBUFX2TS \fifo_from_fft/fifo_cell0/data_out/do_tri[0]  (.Y(fft_data_in[0]), 
	.OE(FE_OFN1142_n585), 
	.A(\fifo_from_fft/fifo_cell0/sr_out[0] ));
   DFFQX1TS \fifo_to_fft/fifo_cell15/hold_token_reg  (.Q(\fifo_to_fft/hold[15] ), 
	.D(\fifo_to_fft/fifo_cell15/N7 ), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell15/hold_token_reg  (.Q(\fifo_to_fir/hold[15] ), 
	.D(\fifo_to_fir/fifo_cell15/N7 ), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/hold_token_reg  (.Q(\fifo_from_fft/hold[15] ), 
	.D(\fifo_from_fft/fifo_cell15/N7 ), 
	.CK(clk__L1_N0));
   TBUFX2TS \router/data_cntl/data_bus_tri[30]  (.Y(data_bus[30]), 
	.OE(FE_OFN994_n521), 
	.A(\router/data_cntl/data_in[30] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[29]  (.Y(data_bus[29]), 
	.OE(FE_OFN997_n521), 
	.A(\router/data_cntl/data_in[29] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[28]  (.Y(data_bus[28]), 
	.OE(FE_OFN997_n521), 
	.A(\router/data_cntl/data_in[28] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[23]  (.Y(data_bus[23]), 
	.OE(FE_OFN1001_n521), 
	.A(\router/data_cntl/data_in[23] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[22]  (.Y(data_bus[22]), 
	.OE(FE_OFN1002_n521), 
	.A(\router/data_cntl/data_in[22] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[21]  (.Y(data_bus[21]), 
	.OE(FE_OFN1001_n521), 
	.A(\router/data_cntl/data_in[21] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[20]  (.Y(data_bus[20]), 
	.OE(FE_OFN1000_n521), 
	.A(\router/data_cntl/data_in[20] ));
   DFFQX1TS \fifo_to_fft/fifo_cell15/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell15/controller/valid_read ), 
	.D(n9519), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell15/controller/valid_read ), 
	.D(n9523), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell15/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell15/controller/valid_read ), 
	.D(n9527), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/iir_write_calc/counter/done_reg  (.Q(\router/iir_write_done ), 
	.D(n6765), 
	.CK(clk__L1_N0));
   DFFTRX2TS \router/addr_calc/from_iir_go_reg  (.RN(\router/data_from_iir ), 
	.QN(\router/addr_calc/N191 ), 
	.Q(n8060), 
	.D(n7607), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell15/reg_ptok/token_reg  (.RN(n4487), 
	.QN(\fifo_from_fft/hang[14] ), 
	.Q(n4598), 
	.D(n4597), 
	.CK(clk__L1_N0));
   TBUFX2TS \router/addr_calc/addr_tri[31]  (.Y(addr[31]), 
	.OE(FE_OFN1218_n8064), 
	.A(n7488));
   TBUFX2TS \router/addr_calc/addr_tri[30]  (.Y(addr[30]), 
	.OE(FE_OFN1218_n8064), 
	.A(FE_OFN1229_router_addr_calc_fft_read_calc_count_30_));
   TBUFX2TS \router/addr_calc/addr_tri[29]  (.Y(addr[29]), 
	.OE(FE_OFN1218_n8064), 
	.A(FE_OFN1234_n7492));
   TBUFX2TS \router/addr_calc/addr_tri[28]  (.Y(addr[28]), 
	.OE(FE_OFN1221_n8064), 
	.A(n7497));
   TBUFX2TS \router/addr_calc/addr_tri[27]  (.Y(addr[27]), 
	.OE(FE_OFN1220_n8064), 
	.A(FE_OFN1237_router_addr_calc_fft_read_calc_count_27_));
   TBUFX2TS \router/addr_calc/addr_tri[26]  (.Y(addr[26]), 
	.OE(FE_OFN1220_n8064), 
	.A(n7502));
   TBUFX2TS \router/addr_calc/addr_tri[25]  (.Y(addr[25]), 
	.OE(FE_OFN1220_n8064), 
	.A(n7506));
   TBUFX2TS \router/addr_calc/addr_tri[24]  (.Y(addr[24]), 
	.OE(FE_OFN1220_n8064), 
	.A(n7511));
   TBUFX2TS \router/addr_calc/addr_tri[23]  (.Y(addr[23]), 
	.OE(FE_OFN857_n7017), 
	.A(FE_OFN1245_router_addr_calc_fft_read_calc_count_23_));
   TBUFX2TS \router/addr_calc/addr_tri[22]  (.Y(addr[22]), 
	.OE(FE_OFN858_n7017), 
	.A(n7516));
   TBUFX2TS \router/addr_calc/addr_tri[21]  (.Y(addr[21]), 
	.OE(FE_OFN858_n7017), 
	.A(n7521));
   TBUFX2TS \router/addr_calc/addr_tri[20]  (.Y(addr[20]), 
	.OE(FE_OFN861_n7017), 
	.A(n7526));
   TBUFX2TS \router/addr_calc/addr_tri[19]  (.Y(addr[19]), 
	.OE(FE_OFN861_n7017), 
	.A(FE_OFN1258_router_addr_calc_fft_read_calc_count_19_));
   TBUFX2TS \router/addr_calc/addr_tri[18]  (.Y(addr[18]), 
	.OE(FE_OFN859_n7017), 
	.A(n7532));
   TBUFX2TS \router/addr_calc/addr_tri[17]  (.Y(addr[17]), 
	.OE(FE_OFN860_n7017), 
	.A(n7536));
   TBUFX2TS \router/addr_calc/addr_tri[16]  (.Y(addr[16]), 
	.OE(FE_OFN860_n7017), 
	.A(FE_OFN1263_router_addr_calc_fft_read_calc_count_16_));
   TBUFX2TS \router/addr_calc/addr_tri[15]  (.Y(addr[15]), 
	.OE(FE_OFN860_n7017), 
	.A(n7541));
   TBUFX2TS \router/addr_calc/addr_tri[14]  (.Y(addr[14]), 
	.OE(FE_OFN861_n7017), 
	.A(n7546));
   TBUFX2TS \router/addr_calc/addr_tri[13]  (.Y(addr[13]), 
	.OE(FE_OFN861_n7017), 
	.A(n7551));
   TBUFX2TS \router/addr_calc/addr_tri[12]  (.Y(addr[12]), 
	.OE(FE_OFN859_n7017), 
	.A(n7556));
   TBUFX2TS \router/addr_calc/addr_tri[11]  (.Y(addr[11]), 
	.OE(FE_OFN859_n7017), 
	.A(n7561));
   TBUFX2TS \router/addr_calc/addr_tri[10]  (.Y(addr[10]), 
	.OE(FE_OFN857_n7017), 
	.A(n7566));
   TBUFX2TS \router/addr_calc/addr_tri[9]  (.Y(addr[9]), 
	.OE(FE_OFN857_n7017), 
	.A(\router/addr_calc/fft_read_calc/count[9] ));
   TBUFX2TS \router/addr_calc/addr_tri[8]  (.Y(addr[8]), 
	.OE(n7017), 
	.A(n7571));
   TBUFX2TS \router/addr_calc/addr_tri[7]  (.Y(addr[7]), 
	.OE(FE_OFN1222_n8064), 
	.A(n7576));
   TBUFX2TS \router/addr_calc/addr_tri[6]  (.Y(addr[6]), 
	.OE(FE_OFN1222_n8064), 
	.A(n7581));
   TBUFX2TS \router/addr_calc/addr_tri[5]  (.Y(addr[5]), 
	.OE(FE_OFN1219_n8064), 
	.A(FE_OFN1273_router_addr_calc_fft_read_calc_count_5_));
   TBUFX2TS \router/addr_calc/addr_tri[4]  (.Y(addr[4]), 
	.OE(FE_OFN1219_n8064), 
	.A(n7587));
   TBUFX2TS \router/addr_calc/addr_tri[3]  (.Y(addr[3]), 
	.OE(n8064), 
	.A(n7591));
   TBUFX2TS \router/addr_calc/addr_tri[2]  (.Y(addr[2]), 
	.OE(n8064), 
	.A(n7596));
   TBUFX2TS \router/addr_calc/addr_tri[1]  (.Y(addr[1]), 
	.OE(FE_OFN1221_n8064), 
	.A(n7602));
   TBUFX2TS \router/addr_calc/addr_tri[0]  (.Y(addr[0]), 
	.OE(FE_OFN1221_n8064), 
	.A(FE_OFN1444_router_addr_calc_fft_read_calc_count_0_));
   TBUFX2TS \router/addr_calc/addr_tri2[31]  (.Y(addr[31]), 
	.OE(FE_OFN1227_n8063), 
	.A(FE_OFN1228_router_addr_calc_fft_write_calc_count_31_));
   TBUFX2TS \router/addr_calc/addr_tri2[30]  (.Y(addr[30]), 
	.OE(n8063), 
	.A(FE_OFN1232_n7368));
   TBUFX2TS \router/addr_calc/addr_tri2[29]  (.Y(addr[29]), 
	.OE(FE_OFN1227_n8063), 
	.A(FE_OFN1233_router_addr_calc_fft_write_calc_count_29_));
   TBUFX2TS \router/addr_calc/addr_tri2[28]  (.Y(addr[28]), 
	.OE(FE_OFN1225_n8063), 
	.A(n7373));
   TBUFX2TS \router/addr_calc/addr_tri2[27]  (.Y(addr[27]), 
	.OE(FE_OFN1223_n8063), 
	.A(FE_OFN1238_router_addr_calc_fft_write_calc_count_27_));
   TBUFX2TS \router/addr_calc/addr_tri2[26]  (.Y(addr[26]), 
	.OE(FE_OFN1224_n8063), 
	.A(n7378));
   TBUFX2TS \router/addr_calc/addr_tri2[25]  (.Y(addr[25]), 
	.OE(FE_OFN1224_n8063), 
	.A(n7382));
   TBUFX2TS \router/addr_calc/addr_tri2[24]  (.Y(addr[24]), 
	.OE(FE_OFN1224_n8063), 
	.A(n7387));
   TBUFX2TS \router/addr_calc/addr_tri2[23]  (.Y(addr[23]), 
	.OE(n7015), 
	.A(FE_OFN1246_router_addr_calc_fft_write_calc_count_23_));
   TBUFX2TS \router/addr_calc/addr_tri2[22]  (.Y(addr[22]), 
	.OE(FE_OFN862_n7015), 
	.A(FE_OFN1249_n7392));
   TBUFX2TS \router/addr_calc/addr_tri2[21]  (.Y(addr[21]), 
	.OE(FE_OFN862_n7015), 
	.A(FE_OFN1252_n7397));
   TBUFX2TS \router/addr_calc/addr_tri2[20]  (.Y(addr[20]), 
	.OE(FE_OFN866_n7015), 
	.A(FE_OFN1255_n7402));
   TBUFX2TS \router/addr_calc/addr_tri2[19]  (.Y(addr[19]), 
	.OE(FE_OFN865_n7015), 
	.A(FE_OFN1259_router_addr_calc_fft_write_calc_count_19_));
   TBUFX2TS \router/addr_calc/addr_tri2[18]  (.Y(addr[18]), 
	.OE(FE_OFN863_n7015), 
	.A(n7408));
   TBUFX2TS \router/addr_calc/addr_tri2[17]  (.Y(addr[17]), 
	.OE(FE_OFN865_n7015), 
	.A(n7412));
   TBUFX2TS \router/addr_calc/addr_tri2[16]  (.Y(addr[16]), 
	.OE(FE_OFN865_n7015), 
	.A(n7417));
   TBUFX2TS \router/addr_calc/addr_tri2[15]  (.Y(addr[15]), 
	.OE(FE_OFN866_n7015), 
	.A(\router/addr_calc/fft_write_calc/count[15] ));
   TBUFX2TS \router/addr_calc/addr_tri2[14]  (.Y(addr[14]), 
	.OE(FE_OFN866_n7015), 
	.A(n7422));
   TBUFX2TS \router/addr_calc/addr_tri2[13]  (.Y(addr[13]), 
	.OE(FE_OFN866_n7015), 
	.A(n7427));
   TBUFX2TS \router/addr_calc/addr_tri2[12]  (.Y(addr[12]), 
	.OE(FE_OFN863_n7015), 
	.A(n7432));
   TBUFX2TS \router/addr_calc/addr_tri2[11]  (.Y(addr[11]), 
	.OE(FE_OFN864_n7015), 
	.A(n7437));
   TBUFX2TS \router/addr_calc/addr_tri2[10]  (.Y(addr[10]), 
	.OE(FE_OFN864_n7015), 
	.A(n7442));
   TBUFX2TS \router/addr_calc/addr_tri2[9]  (.Y(addr[9]), 
	.OE(FE_OFN864_n7015), 
	.A(FE_OFN1268_router_addr_calc_fft_write_calc_count_9_));
   TBUFX2TS \router/addr_calc/addr_tri2[8]  (.Y(addr[8]), 
	.OE(FE_OFN864_n7015), 
	.A(n7447));
   TBUFX2TS \router/addr_calc/addr_tri2[7]  (.Y(addr[7]), 
	.OE(FE_OFN1226_n8063), 
	.A(n7452));
   TBUFX2TS \router/addr_calc/addr_tri2[6]  (.Y(addr[6]), 
	.OE(FE_OFN1227_n8063), 
	.A(n7457));
   TBUFX2TS \router/addr_calc/addr_tri2[5]  (.Y(addr[5]), 
	.OE(FE_OFN1223_n8063), 
	.A(n7463));
   TBUFX2TS \router/addr_calc/addr_tri2[4]  (.Y(addr[4]), 
	.OE(FE_OFN1226_n8063), 
	.A(n7468));
   TBUFX2TS \router/addr_calc/addr_tri2[3]  (.Y(addr[3]), 
	.OE(FE_OFN1225_n8063), 
	.A(n7472));
   TBUFX2TS \router/addr_calc/addr_tri2[2]  (.Y(addr[2]), 
	.OE(FE_OFN1225_n8063), 
	.A(n7477));
   TBUFX2TS \router/addr_calc/addr_tri2[1]  (.Y(addr[1]), 
	.OE(FE_OFN1224_n8063), 
	.A(n7483));
   TBUFX2TS \router/addr_calc/addr_tri2[0]  (.Y(addr[0]), 
	.OE(FE_OFN1226_n8063), 
	.A(FE_OFN1443_router_addr_calc_fft_write_calc_count_0_));
   TBUFX2TS \router/addr_calc/addr_tri3[31]  (.Y(addr[31]), 
	.OE(n8062), 
	.A(n7250));
   TBUFX2TS \router/addr_calc/addr_tri3[30]  (.Y(addr[30]), 
	.OE(n8062), 
	.A(FE_OFN1230_router_addr_calc_fir_read_calc_count_30_));
   TBUFX2TS \router/addr_calc/addr_tri3[29]  (.Y(addr[29]), 
	.OE(n8062), 
	.A(FE_OFN1235_n7254));
   TBUFX2TS \router/addr_calc/addr_tri3[28]  (.Y(addr[28]), 
	.OE(FE_OFN1209_n8062), 
	.A(FE_OFN1236_n7259));
   TBUFX2TS \router/addr_calc/addr_tri3[27]  (.Y(addr[27]), 
	.OE(FE_OFN1210_n8062), 
	.A(FE_OFN1239_router_addr_calc_fir_read_calc_count_27_));
   TBUFX2TS \router/addr_calc/addr_tri3[26]  (.Y(addr[26]), 
	.OE(FE_OFN1211_n8062), 
	.A(FE_OFN1241_n7264));
   TBUFX2TS \router/addr_calc/addr_tri3[25]  (.Y(addr[25]), 
	.OE(FE_OFN1211_n8062), 
	.A(FE_OFN1242_n7268));
   TBUFX2TS \router/addr_calc/addr_tri3[24]  (.Y(addr[24]), 
	.OE(FE_OFN1211_n8062), 
	.A(FE_OFN1243_n7273));
   TBUFX2TS \router/addr_calc/addr_tri3[23]  (.Y(addr[23]), 
	.OE(FE_OFN850_n7016), 
	.A(FE_OFN1247_router_addr_calc_fir_read_calc_count_23_));
   TBUFX2TS \router/addr_calc/addr_tri3[22]  (.Y(addr[22]), 
	.OE(FE_OFN849_n7016), 
	.A(FE_OFN1250_n7278));
   TBUFX2TS \router/addr_calc/addr_tri3[21]  (.Y(addr[21]), 
	.OE(FE_OFN850_n7016), 
	.A(FE_OFN1253_n7283));
   TBUFX2TS \router/addr_calc/addr_tri3[20]  (.Y(addr[20]), 
	.OE(FE_OFN851_n7016), 
	.A(FE_OFN1256_n7288));
   TBUFX2TS \router/addr_calc/addr_tri3[19]  (.Y(addr[19]), 
	.OE(FE_OFN852_n7016), 
	.A(FE_OFN1260_router_addr_calc_fir_read_calc_count_19_));
   TBUFX2TS \router/addr_calc/addr_tri3[18]  (.Y(addr[18]), 
	.OE(FE_OFN849_n7016), 
	.A(n7294));
   TBUFX2TS \router/addr_calc/addr_tri3[17]  (.Y(addr[17]), 
	.OE(FE_OFN852_n7016), 
	.A(FE_OFN1262_n7298));
   TBUFX2TS \router/addr_calc/addr_tri3[16]  (.Y(addr[16]), 
	.OE(FE_OFN852_n7016), 
	.A(FE_OFN1265_n7303));
   TBUFX2TS \router/addr_calc/addr_tri3[15]  (.Y(addr[15]), 
	.OE(FE_OFN852_n7016), 
	.A(\router/addr_calc/fir_read_calc/count[15] ));
   TBUFX2TS \router/addr_calc/addr_tri3[14]  (.Y(addr[14]), 
	.OE(FE_OFN851_n7016), 
	.A(FE_OFN1277_n7308));
   TBUFX2TS \router/addr_calc/addr_tri3[13]  (.Y(addr[13]), 
	.OE(FE_OFN851_n7016), 
	.A(n7313));
   TBUFX2TS \router/addr_calc/addr_tri3[12]  (.Y(addr[12]), 
	.OE(FE_OFN850_n7016), 
	.A(n7318));
   TBUFX2TS \router/addr_calc/addr_tri3[11]  (.Y(addr[11]), 
	.OE(FE_OFN849_n7016), 
	.A(n7323));
   TBUFX2TS \router/addr_calc/addr_tri3[10]  (.Y(addr[10]), 
	.OE(n7016), 
	.A(FE_OFN1279_n7328));
   TBUFX2TS \router/addr_calc/addr_tri3[9]  (.Y(addr[9]), 
	.OE(n7016), 
	.A(FE_OFN1269_router_addr_calc_fir_read_calc_count_9_));
   TBUFX2TS \router/addr_calc/addr_tri3[8]  (.Y(addr[8]), 
	.OE(n7016), 
	.A(FE_OFN1278_n7333));
   TBUFX2TS \router/addr_calc/addr_tri3[7]  (.Y(addr[7]), 
	.OE(FE_OFN1210_n8062), 
	.A(n7338));
   TBUFX2TS \router/addr_calc/addr_tri3[6]  (.Y(addr[6]), 
	.OE(FE_OFN1210_n8062), 
	.A(n7343));
   TBUFX2TS \router/addr_calc/addr_tri3[5]  (.Y(addr[5]), 
	.OE(FE_OFN1208_n8062), 
	.A(FE_OFN1824_router_addr_calc_fir_read_calc_count_5_));
   TBUFX2TS \router/addr_calc/addr_tri3[4]  (.Y(addr[4]), 
	.OE(FE_OFN1211_n8062), 
	.A(n7349));
   TBUFX2TS \router/addr_calc/addr_tri3[3]  (.Y(addr[3]), 
	.OE(FE_OFN1208_n8062), 
	.A(FE_OFN1275_n7353));
   TBUFX2TS \router/addr_calc/addr_tri3[2]  (.Y(addr[2]), 
	.OE(FE_OFN1208_n8062), 
	.A(FE_OFN1274_n7358));
   TBUFX2TS \router/addr_calc/addr_tri3[1]  (.Y(addr[1]), 
	.OE(FE_OFN1209_n8062), 
	.A(n7364));
   TBUFX2TS \router/addr_calc/addr_tri3[0]  (.Y(addr[0]), 
	.OE(FE_OFN1210_n8062), 
	.A(FE_OFN1446_router_addr_calc_fir_read_calc_count_0_));
   TBUFX2TS \router/addr_calc/addr_tri4[31]  (.Y(addr[31]), 
	.OE(n8061), 
	.A(n7119));
   TBUFX2TS \router/addr_calc/addr_tri4[30]  (.Y(addr[30]), 
	.OE(FE_OFN1213_n8061), 
	.A(FE_OFN1231_router_addr_calc_fir_write_calc_count_30_));
   TBUFX2TS \router/addr_calc/addr_tri4[29]  (.Y(addr[29]), 
	.OE(n8061), 
	.A(n7124));
   TBUFX2TS \router/addr_calc/addr_tri4[28]  (.Y(addr[28]), 
	.OE(FE_OFN1213_n8061), 
	.A(n7130));
   TBUFX2TS \router/addr_calc/addr_tri4[27]  (.Y(addr[27]), 
	.OE(FE_OFN1215_n8061), 
	.A(FE_OFN1240_router_addr_calc_fir_write_calc_count_27_));
   TBUFX2TS \router/addr_calc/addr_tri4[26]  (.Y(addr[26]), 
	.OE(FE_OFN1213_n8061), 
	.A(n7136));
   TBUFX2TS \router/addr_calc/addr_tri4[25]  (.Y(addr[25]), 
	.OE(FE_OFN1216_n8061), 
	.A(n7141));
   TBUFX2TS \router/addr_calc/addr_tri4[24]  (.Y(addr[24]), 
	.OE(FE_OFN1216_n8061), 
	.A(n7147));
   TBUFX2TS \router/addr_calc/addr_tri4[23]  (.Y(addr[23]), 
	.OE(n7018), 
	.A(FE_OFN1248_router_addr_calc_fir_write_calc_count_23_));
   TBUFX2TS \router/addr_calc/addr_tri4[22]  (.Y(addr[22]), 
	.OE(FE_OFN853_n7018), 
	.A(FE_OFN1251_n7153));
   TBUFX2TS \router/addr_calc/addr_tri4[21]  (.Y(addr[21]), 
	.OE(FE_OFN853_n7018), 
	.A(FE_OFN1254_n7159));
   TBUFX2TS \router/addr_calc/addr_tri4[20]  (.Y(addr[20]), 
	.OE(FE_OFN855_n7018), 
	.A(FE_OFN1257_n7165));
   TBUFX2TS \router/addr_calc/addr_tri4[19]  (.Y(addr[19]), 
	.OE(FE_OFN855_n7018), 
	.A(FE_OFN1261_router_addr_calc_fir_write_calc_count_19_));
   TBUFX2TS \router/addr_calc/addr_tri4[18]  (.Y(addr[18]), 
	.OE(FE_OFN855_n7018), 
	.A(n7172));
   TBUFX2TS \router/addr_calc/addr_tri4[17]  (.Y(addr[17]), 
	.OE(FE_OFN854_n7018), 
	.A(n7177));
   TBUFX2TS \router/addr_calc/addr_tri4[16]  (.Y(addr[16]), 
	.OE(FE_OFN856_n7018), 
	.A(FE_OFN1264_router_addr_calc_fir_write_calc_count_16_));
   TBUFX2TS \router/addr_calc/addr_tri4[15]  (.Y(addr[15]), 
	.OE(FE_OFN856_n7018), 
	.A(n7183));
   TBUFX2TS \router/addr_calc/addr_tri4[14]  (.Y(addr[14]), 
	.OE(FE_OFN856_n7018), 
	.A(n7189));
   TBUFX2TS \router/addr_calc/addr_tri4[13]  (.Y(addr[13]), 
	.OE(FE_OFN856_n7018), 
	.A(n7195));
   TBUFX2TS \router/addr_calc/addr_tri4[12]  (.Y(addr[12]), 
	.OE(FE_OFN854_n7018), 
	.A(n7201));
   TBUFX2TS \router/addr_calc/addr_tri4[11]  (.Y(addr[11]), 
	.OE(FE_OFN854_n7018), 
	.A(n7205));
   TBUFX2TS \router/addr_calc/addr_tri4[10]  (.Y(addr[10]), 
	.OE(FE_OFN854_n7018), 
	.A(n7209));
   TBUFX2TS \router/addr_calc/addr_tri4[9]  (.Y(addr[9]), 
	.OE(n7018), 
	.A(FE_OFN1266_router_addr_calc_fir_write_calc_count_9_));
   TBUFX2TS \router/addr_calc/addr_tri4[8]  (.Y(addr[8]), 
	.OE(n7018), 
	.A(n7214));
   TBUFX2TS \router/addr_calc/addr_tri4[7]  (.Y(addr[7]), 
	.OE(FE_OFN1216_n8061), 
	.A(n7219));
   TBUFX2TS \router/addr_calc/addr_tri4[6]  (.Y(addr[6]), 
	.OE(FE_OFN1215_n8061), 
	.A(n7224));
   TBUFX2TS \router/addr_calc/addr_tri4[5]  (.Y(addr[5]), 
	.OE(FE_OFN1214_n8061), 
	.A(FE_OFN1272_router_addr_calc_fir_write_calc_count_5_));
   TBUFX2TS \router/addr_calc/addr_tri4[4]  (.Y(addr[4]), 
	.OE(FE_OFN1214_n8061), 
	.A(n7230));
   TBUFX2TS \router/addr_calc/addr_tri4[3]  (.Y(addr[3]), 
	.OE(FE_OFN1212_n8061), 
	.A(n7234));
   TBUFX2TS \router/addr_calc/addr_tri4[2]  (.Y(addr[2]), 
	.OE(FE_OFN1214_n8061), 
	.A(n7239));
   TBUFX2TS \router/addr_calc/addr_tri4[1]  (.Y(addr[1]), 
	.OE(FE_OFN1215_n8061), 
	.A(n7245));
   TBUFX2TS \router/addr_calc/addr_tri4[0]  (.Y(addr[0]), 
	.OE(FE_OFN1212_n8061), 
	.A(FE_OFN1445_router_addr_calc_fir_write_calc_count_0_));
   TBUFX2TS \router/addr_calc/addr_tri5[31]  (.Y(addr[31]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[31] ));
   TBUFX2TS \router/addr_calc/addr_tri5[30]  (.Y(addr[30]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[30] ));
   TBUFX2TS \router/addr_calc/addr_tri5[29]  (.Y(addr[29]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[29] ));
   TBUFX2TS \router/addr_calc/addr_tri5[28]  (.Y(addr[28]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[28] ));
   TBUFX2TS \router/addr_calc/addr_tri5[27]  (.Y(addr[27]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[27] ));
   TBUFX2TS \router/addr_calc/addr_tri5[26]  (.Y(addr[26]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[26] ));
   TBUFX2TS \router/addr_calc/addr_tri5[25]  (.Y(addr[25]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[25] ));
   TBUFX2TS \router/addr_calc/addr_tri5[24]  (.Y(addr[24]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[24] ));
   TBUFX2TS \router/addr_calc/addr_tri5[23]  (.Y(addr[23]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[23] ));
   TBUFX2TS \router/addr_calc/addr_tri5[22]  (.Y(addr[22]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[22] ));
   TBUFX2TS \router/addr_calc/addr_tri5[21]  (.Y(addr[21]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[21] ));
   TBUFX2TS \router/addr_calc/addr_tri5[20]  (.Y(addr[20]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[20] ));
   TBUFX2TS \router/addr_calc/addr_tri5[19]  (.Y(addr[19]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[19] ));
   TBUFX2TS \router/addr_calc/addr_tri5[18]  (.Y(addr[18]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[18] ));
   TBUFX2TS \router/addr_calc/addr_tri5[17]  (.Y(addr[17]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[17] ));
   TBUFX2TS \router/addr_calc/addr_tri5[16]  (.Y(addr[16]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[16] ));
   TBUFX2TS \router/addr_calc/addr_tri5[15]  (.Y(addr[15]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[15] ));
   TBUFX2TS \router/addr_calc/addr_tri5[14]  (.Y(addr[14]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[14] ));
   TBUFX2TS \router/addr_calc/addr_tri5[13]  (.Y(addr[13]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[13] ));
   TBUFX2TS \router/addr_calc/addr_tri5[12]  (.Y(addr[12]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[12] ));
   TBUFX2TS \router/addr_calc/addr_tri5[11]  (.Y(addr[11]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[11] ));
   TBUFX2TS \router/addr_calc/addr_tri5[10]  (.Y(addr[10]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[10] ));
   TBUFX2TS \router/addr_calc/addr_tri5[9]  (.Y(addr[9]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[9] ));
   TBUFX2TS \router/addr_calc/addr_tri5[8]  (.Y(addr[8]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[8] ));
   TBUFX2TS \router/addr_calc/addr_tri5[7]  (.Y(addr[7]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[7] ));
   TBUFX2TS \router/addr_calc/addr_tri5[6]  (.Y(addr[6]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[6] ));
   TBUFX2TS \router/addr_calc/addr_tri5[5]  (.Y(addr[5]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[5] ));
   TBUFX2TS \router/addr_calc/addr_tri5[4]  (.Y(addr[4]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[4] ));
   TBUFX2TS \router/addr_calc/addr_tri5[3]  (.Y(addr[3]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[3] ));
   TBUFX2TS \router/addr_calc/addr_tri5[2]  (.Y(addr[2]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[2] ));
   TBUFX2TS \router/addr_calc/addr_tri5[1]  (.Y(addr[1]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[1] ));
   TBUFX2TS \router/addr_calc/addr_tri5[0]  (.Y(addr[0]), 
	.OE(1'b0), 
	.A(\router/addr_calc/iir_read_calc/count[0] ));
   TBUFX2TS \router/addr_calc/addr_tri6[31]  (.Y(addr[31]), 
	.OE(FE_OFN1305_n8060), 
	.A(n7199));
   TBUFX2TS \router/addr_calc/addr_tri6[29]  (.Y(addr[29]), 
	.OE(FE_OFN1305_n8060), 
	.A(n7193));
   TBUFX2TS \router/addr_calc/addr_tri6[28]  (.Y(addr[28]), 
	.OE(FE_OFN1302_n8060), 
	.A(n7187));
   TBUFX2TS \router/addr_calc/addr_tri6[27]  (.Y(addr[27]), 
	.OE(FE_OFN1302_n8060), 
	.A(\router/addr_calc/iir_write_calc/count[27] ));
   TBUFX2TS \router/addr_calc/addr_tri6[26]  (.Y(addr[26]), 
	.OE(FE_OFN1301_n8060), 
	.A(n7181));
   TBUFX2TS \router/addr_calc/addr_tri6[25]  (.Y(addr[25]), 
	.OE(FE_OFN1301_n8060), 
	.A(n7174));
   TBUFX2TS \router/addr_calc/addr_tri6[24]  (.Y(addr[24]), 
	.OE(FE_OFN1301_n8060), 
	.A(n7168));
   TBUFX2TS \router/addr_calc/addr_tri6[23]  (.Y(addr[23]), 
	.OE(FE_OFN1007_n137), 
	.A(FE_OFN1244_router_addr_calc_iir_write_calc_count_23_));
   TBUFX2TS \router/addr_calc/addr_tri6[22]  (.Y(addr[22]), 
	.OE(FE_OFN1007_n137), 
	.A(n7162));
   TBUFX2TS \router/addr_calc/addr_tri6[21]  (.Y(addr[21]), 
	.OE(FE_OFN1007_n137), 
	.A(n7156));
   TBUFX2TS \router/addr_calc/addr_tri6[20]  (.Y(addr[20]), 
	.OE(FE_OFN1005_n137), 
	.A(n7150));
   TBUFX2TS \router/addr_calc/addr_tri6[19]  (.Y(addr[19]), 
	.OE(FE_OFN1008_n137), 
	.A(\router/addr_calc/iir_write_calc/count[19] ));
   TBUFX2TS \router/addr_calc/addr_tri6[18]  (.Y(addr[18]), 
	.OE(FE_OFN1006_n137), 
	.A(n7145));
   TBUFX2TS \router/addr_calc/addr_tri6[17]  (.Y(addr[17]), 
	.OE(FE_OFN1008_n137), 
	.A(n7138));
   TBUFX2TS \router/addr_calc/addr_tri6[16]  (.Y(addr[16]), 
	.OE(FE_OFN1008_n137), 
	.A(\router/addr_calc/iir_write_calc/count[16] ));
   TBUFX2TS \router/addr_calc/addr_tri6[15]  (.Y(addr[15]), 
	.OE(FE_OFN1005_n137), 
	.A(n7132));
   TBUFX2TS \router/addr_calc/addr_tri6[14]  (.Y(addr[14]), 
	.OE(FE_OFN1008_n137), 
	.A(n7126));
   TBUFX2TS \router/addr_calc/addr_tri6[13]  (.Y(addr[13]), 
	.OE(FE_OFN1005_n137), 
	.A(n7121));
   TBUFX2TS \router/addr_calc/addr_tri6[12]  (.Y(addr[12]), 
	.OE(FE_OFN1006_n137), 
	.A(n7115));
   TBUFX2TS \router/addr_calc/addr_tri6[11]  (.Y(addr[11]), 
	.OE(FE_OFN1006_n137), 
	.A(n7109));
   TBUFX2TS \router/addr_calc/addr_tri6[10]  (.Y(addr[10]), 
	.OE(FE_OFN1004_n137), 
	.A(n7104));
   TBUFX2TS \router/addr_calc/addr_tri6[9]  (.Y(addr[9]), 
	.OE(n137), 
	.A(FE_OFN1280_router_addr_calc_iir_write_calc_count_9_));
   TBUFX2TS \router/addr_calc/addr_tri6[8]  (.Y(addr[8]), 
	.OE(FE_OFN1004_n137), 
	.A(n7098));
   TBUFX2TS \router/addr_calc/addr_tri6[7]  (.Y(addr[7]), 
	.OE(FE_OFN1303_n8060), 
	.A(n7092));
   TBUFX2TS \router/addr_calc/addr_tri6[6]  (.Y(addr[6]), 
	.OE(FE_OFN1303_n8060), 
	.A(n7089));
   TBUFX2TS \router/addr_calc/addr_tri6[5]  (.Y(addr[5]), 
	.OE(FE_OFN1304_n8060), 
	.A(\router/addr_calc/iir_write_calc/count[5] ));
   TBUFX2TS \router/addr_calc/addr_tri6[4]  (.Y(addr[4]), 
	.OE(FE_OFN1305_n8060), 
	.A(n7096));
   TBUFX2TS \router/addr_calc/addr_tri6[3]  (.Y(addr[3]), 
	.OE(FE_OFN1304_n8060), 
	.A(n7101));
   TBUFX2TS \router/addr_calc/addr_tri6[1]  (.Y(addr[1]), 
	.OE(n8060), 
	.A(n7113));
   TBUFX2TS \router/addr_calc/addr_tri6[0]  (.Y(addr[0]), 
	.OE(FE_OFN1303_n8060), 
	.A(FE_OFN1442_router_addr_calc_iir_write_calc_count_0_));
   DFFQX1TS \fifo_from_fir/fifo_cell15/hold_token_reg  (.Q(\fifo_from_fir/hold[15] ), 
	.D(\fifo_from_fir/fifo_cell15/N7 ), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/ram_write_reg  (.Q(\router/ram_write_enable_reg ), 
	.D(n6763), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/iir_full_flag_reg  (.Q(\router/data_cntl/N151 ), 
	.D(n5461), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell13/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell13/reg_gtok/token ), 
	.D(n5475), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell14/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell14/reg_gtok/token ), 
	.D(n5472), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell13/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell13/reg_gtok/token ), 
	.D(n5527), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell14/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell14/reg_gtok/token ), 
	.D(n5524), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell14/reg_gtok/token ), 
	.D(n6746), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell14/reg_gtok/token ), 
	.D(n6217), 
	.CK(clk__L1_N0));
   TBUFX2TS \router/data_cntl/data_bus_tri[27]  (.Y(data_bus[27]), 
	.OE(FE_OFN994_n521), 
	.A(\router/data_cntl/data_in[27] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[26]  (.Y(data_bus[26]), 
	.OE(FE_OFN998_n521), 
	.A(\router/data_cntl/data_in[26] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[25]  (.Y(data_bus[25]), 
	.OE(n521), 
	.A(\router/data_cntl/data_in[25] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[24]  (.Y(data_bus[24]), 
	.OE(n521), 
	.A(\router/data_cntl/data_in[24] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[19]  (.Y(data_bus[19]), 
	.OE(FE_OFN998_n521), 
	.A(\router/data_cntl/data_in[19] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[18]  (.Y(data_bus[18]), 
	.OE(FE_OFN999_n521), 
	.A(\router/data_cntl/data_in[18] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[17]  (.Y(data_bus[17]), 
	.OE(FE_OFN999_n521), 
	.A(\router/data_cntl/data_in[17] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[16]  (.Y(data_bus[16]), 
	.OE(FE_OFN997_n521), 
	.A(\router/data_cntl/data_in[16] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[15]  (.Y(data_bus[15]), 
	.OE(FE_OFN1002_n521), 
	.A(\router/data_cntl/data_in[15] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[14]  (.Y(data_bus[14]), 
	.OE(FE_OFN1000_n521), 
	.A(\router/data_cntl/data_in[14] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[13]  (.Y(data_bus[13]), 
	.OE(FE_OFN1003_n521), 
	.A(\router/data_cntl/data_in[13] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[12]  (.Y(data_bus[12]), 
	.OE(FE_OFN1000_n521), 
	.A(\router/data_cntl/data_in[12] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[11]  (.Y(data_bus[11]), 
	.OE(FE_OFN1003_n521), 
	.A(\router/data_cntl/data_in[11] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[10]  (.Y(data_bus[10]), 
	.OE(FE_OFN1001_n521), 
	.A(\router/data_cntl/data_in[10] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[9]  (.Y(data_bus[9]), 
	.OE(FE_OFN1003_n521), 
	.A(\router/data_cntl/data_in[9] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[8]  (.Y(data_bus[8]), 
	.OE(FE_OFN1002_n521), 
	.A(\router/data_cntl/data_in[8] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[7]  (.Y(data_bus[7]), 
	.OE(FE_OFN994_n521), 
	.A(\router/data_cntl/data_in[7] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[6]  (.Y(data_bus[6]), 
	.OE(FE_OFN996_n521), 
	.A(\router/data_cntl/data_in[6] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[5]  (.Y(data_bus[5]), 
	.OE(n521), 
	.A(\router/data_cntl/data_in[5] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[4]  (.Y(data_bus[4]), 
	.OE(FE_OFN995_n521), 
	.A(\router/data_cntl/data_in[4] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[3]  (.Y(data_bus[3]), 
	.OE(FE_OFN998_n521), 
	.A(\router/data_cntl/data_in[3] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[2]  (.Y(data_bus[2]), 
	.OE(FE_OFN996_n521), 
	.A(\router/data_cntl/data_in[2] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[1]  (.Y(data_bus[1]), 
	.OE(FE_OFN995_n521), 
	.A(\router/data_cntl/data_in[1] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[0]  (.Y(data_bus[0]), 
	.OE(FE_OFN999_n521), 
	.A(\router/data_cntl/data_in[0] ));
   TBUFX2TS \router/data_cntl/data_bus_tri[31]  (.Y(data_bus[31]), 
	.OE(FE_OFN995_n521), 
	.A(\router/data_cntl/data_in[31] ));
   DFFQX1TS \fifo_to_fir/fifo_cell0/reg_ptok/token_reg  (.Q(\fifo_to_fir/tok_xnor_put ), 
	.D(n5570), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell0/reg_ptok/token_reg  (.Q(\fifo_to_fft/tok_xnor_put ), 
	.D(n5518), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/fft_full_flag_reg  (.Q(\router/data_cntl/fft_full_flag ), 
	.D(n5460), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell14/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell14/controller/valid_read ), 
	.D(n9519), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell14/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell14/controller/valid_read ), 
	.D(n9527), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell15/controller/valid_read ), 
	.D(n9516), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell15/reg_ptok/token_reg  (.RN(n4673), 
	.QN(\fifo_from_fir/hang[14] ), 
	.Q(n4784), 
	.D(n4783), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell14/reg_ptok/token_reg  (.RN(n3878), 
	.QN(\fifo_to_fft/hang[13] ), 
	.Q(n3964), 
	.D(n3963), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell14/reg_ptok/token_reg  (.RN(n4053), 
	.QN(\fifo_to_fir/hang[13] ), 
	.Q(n4139), 
	.D(n4138), 
	.CK(clk__L1_N0));
   TBUFX2TS \router/addr_calc/addr_tri6[30]  (.Y(addr[30]), 
	.OE(n8060), 
	.A(\router/addr_calc/iir_write_calc/count[30] ));
   TBUFX2TS \router/addr_calc/addr_tri6[2]  (.Y(addr[2]), 
	.OE(FE_OFN1304_n8060), 
	.A(FE_OFN1825_n7107));
   DFFQX1TS \router/pla_top/iir_enable_reg  (.Q(iir_enable), 
	.D(n6764), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell11/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell11/reg_gtok/token ), 
	.D(n5481), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell12/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell12/reg_gtok/token ), 
	.D(n5478), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell11/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell11/reg_gtok/token ), 
	.D(n5533), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell12/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell12/reg_gtok/token ), 
	.D(n5530), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell13/reg_gtok/token ), 
	.D(n6218), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/iir_get_req_reg  (.Q(\router/iir_get_req_reg ), 
	.D(n6762), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/reg_ptok/token_reg  (.Q(\fifo_from_fft/tok_xnor_put ), 
	.D(n5419), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell13/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell13/controller/valid_read ), 
	.D(n9519), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell14/controller/valid_read ), 
	.D(n9523), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell13/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell13/controller/valid_read ), 
	.D(n9527), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell14/reg_ptok/token_reg  (.RN(n4671), 
	.QN(\fifo_from_fir/hang[13] ), 
	.Q(n4787), 
	.D(n4786), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell12/reg_ptok/token_reg  (.RN(n3874), 
	.QN(\fifo_to_fft/hang[11] ), 
	.Q(n3970), 
	.D(n3969), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell13/reg_ptok/token_reg  (.RN(n3876), 
	.QN(\fifo_to_fft/hang[12] ), 
	.Q(n3967), 
	.D(n3966), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell12/reg_ptok/token_reg  (.RN(n4049), 
	.QN(\fifo_to_fir/hang[11] ), 
	.Q(n4145), 
	.D(n4144), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell13/reg_ptok/token_reg  (.RN(n4051), 
	.QN(\fifo_to_fir/hang[12] ), 
	.Q(n4142), 
	.D(n4141), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell14/reg_ptok/token_reg  (.RN(n4485), 
	.QN(\fifo_from_fft/hang[13] ), 
	.Q(n4601), 
	.D(n4600), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/ram_read_reg  (.Q(\router/ram_read_enable_reg ), 
	.D(n6233), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell13/reg_gtok/token ), 
	.D(n6747), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/reg_ptok/token_reg  (.Q(\fifo_from_fir/tok_xnor_put ), 
	.D(n5384), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell11/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell11/controller/valid_read ), 
	.D(n9518), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell12/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell12/controller/valid_read ), 
	.D(n9527), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell11/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell11/controller/valid_read ), 
	.D(n9526), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell12/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell12/controller/valid_read ), 
	.D(n9526), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell14/controller/valid_read ), 
	.D(n9529), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell11/reg_ptok/token_reg  (.RN(n3872), 
	.QN(\fifo_to_fft/hang[10] ), 
	.Q(n3973), 
	.D(n3972), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell11/reg_ptok/token_reg  (.RN(n4047), 
	.QN(\fifo_to_fir/hang[10] ), 
	.Q(n4148), 
	.D(n4147), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell13/reg_ptok/token_reg  (.RN(n4483), 
	.QN(\fifo_from_fft/hang[12] ), 
	.Q(n4604), 
	.D(n4603), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell9/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell9/reg_gtok/token ), 
	.D(n5487), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell10/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell10/reg_gtok/token ), 
	.D(n5484), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell9/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell9/reg_gtok/token ), 
	.D(n5539), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell10/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell10/reg_gtok/token ), 
	.D(n5536), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell12/reg_gtok/token ), 
	.D(n6748), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell12/reg_gtok/token ), 
	.D(n6219), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell10/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell10/controller/valid_read ), 
	.D(n9518), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell13/controller/valid_read ), 
	.D(n9523), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell10/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell10/controller/valid_read ), 
	.D(n9516), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell13/controller/valid_read ), 
	.D(n9531), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell13/reg_ptok/token_reg  (.RN(n4669), 
	.QN(\fifo_from_fir/hang[12] ), 
	.Q(n4790), 
	.D(n4789), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell9/reg_ptok/token_reg  (.RN(n3868), 
	.QN(\fifo_to_fft/hang[8] ), 
	.Q(n3979), 
	.D(n3978), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell10/reg_ptok/token_reg  (.RN(n3870), 
	.QN(\fifo_to_fft/hang[9] ), 
	.Q(n3976), 
	.D(n3975), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell9/reg_ptok/token_reg  (.RN(n4043), 
	.QN(\fifo_to_fir/hang[8] ), 
	.Q(n4154), 
	.D(n4153), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell10/reg_ptok/token_reg  (.RN(n4045), 
	.QN(\fifo_to_fir/hang[9] ), 
	.Q(n4151), 
	.D(n4150), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell7/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell7/reg_gtok/token ), 
	.D(n5493), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell8/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell8/reg_gtok/token ), 
	.D(n5490), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell7/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell7/reg_gtok/token ), 
	.D(n5545), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell8/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell8/reg_gtok/token ), 
	.D(n5542), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell11/reg_gtok/token ), 
	.D(n6220), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell8/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell8/controller/valid_read ), 
	.D(n9518), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell9/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell9/controller/valid_read ), 
	.D(n9518), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell12/controller/valid_read ), 
	.D(n9523), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell8/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell8/controller/valid_read ), 
	.D(n9526), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell9/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell9/controller/valid_read ), 
	.D(n9526), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell12/controller/valid_read ), 
	.D(n9531), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell12/reg_ptok/token_reg  (.RN(n4667), 
	.QN(\fifo_from_fir/hang[11] ), 
	.Q(n4793), 
	.D(n4792), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell12/reg_ptok/token_reg  (.RN(n4481), 
	.QN(\fifo_from_fft/hang[11] ), 
	.Q(n4607), 
	.D(n4606), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell8/reg_ptok/token_reg  (.RN(n3866), 
	.QN(\fifo_to_fft/hang[7] ), 
	.Q(n3982), 
	.D(n3981), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell8/reg_ptok/token_reg  (.RN(n4041), 
	.QN(\fifo_to_fir/hang[7] ), 
	.Q(n4157), 
	.D(n4156), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell6/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell6/reg_gtok/token ), 
	.D(n5496), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell6/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell6/reg_gtok/token ), 
	.D(n5548), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell11/reg_gtok/token ), 
	.D(n6749), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell7/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell7/controller/valid_read ), 
	.D(n9517), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell11/controller/valid_read ), 
	.D(n9522), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell7/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell7/controller/valid_read ), 
	.D(n9525), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell11/reg_ptok/token_reg  (.RN(n4665), 
	.QN(\fifo_from_fir/hang[10] ), 
	.Q(n4796), 
	.D(n4795), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell6/reg_ptok/token_reg  (.RN(n3862), 
	.QN(\fifo_to_fft/hang[5] ), 
	.Q(n3988), 
	.D(n3987), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell7/reg_ptok/token_reg  (.RN(n3864), 
	.QN(\fifo_to_fft/hang[6] ), 
	.Q(n3985), 
	.D(n3984), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell6/reg_ptok/token_reg  (.RN(n4037), 
	.QN(\fifo_to_fir/hang[5] ), 
	.Q(n4163), 
	.D(n4162), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell7/reg_ptok/token_reg  (.RN(n4039), 
	.QN(\fifo_to_fir/hang[6] ), 
	.Q(n4160), 
	.D(n4159), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell11/reg_ptok/token_reg  (.RN(n4479), 
	.QN(\fifo_from_fft/hang[10] ), 
	.Q(n4610), 
	.D(n4609), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell5/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell5/reg_gtok/token ), 
	.D(n5499), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell5/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell5/reg_gtok/token ), 
	.D(n5551), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell10/reg_gtok/token ), 
	.D(n6750), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell10/reg_gtok/token ), 
	.D(n6221), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell5/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell5/controller/valid_read ), 
	.D(n9517), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell6/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell6/controller/valid_read ), 
	.D(n9517), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell5/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell5/controller/valid_read ), 
	.D(n9525), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell6/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell6/controller/valid_read ), 
	.D(n9525), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell11/controller/valid_read ), 
	.D(n9529), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell10/reg_ptok/token_reg  (.RN(n4663), 
	.QN(\fifo_from_fir/hang[9] ), 
	.Q(n4799), 
	.D(n4798), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell5/reg_ptok/token_reg  (.RN(n3860), 
	.QN(\fifo_to_fft/hang[4] ), 
	.Q(n3991), 
	.D(n3990), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell5/reg_ptok/token_reg  (.RN(n4035), 
	.QN(\fifo_to_fir/hang[4] ), 
	.Q(n4166), 
	.D(n4165), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell10/reg_ptok/token_reg  (.RN(n4477), 
	.QN(\fifo_from_fft/hang[9] ), 
	.Q(n4613), 
	.D(n4612), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell3/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell3/reg_gtok/token ), 
	.D(n5505), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell4/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell4/reg_gtok/token ), 
	.D(n5502), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell3/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell3/reg_gtok/token ), 
	.D(n5557), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell4/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell4/reg_gtok/token ), 
	.D(n5554), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell9/reg_gtok/token ), 
	.D(n6751), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell9/reg_gtok/token ), 
	.D(n6222), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell4/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell4/controller/valid_read ), 
	.D(n9517), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell10/controller/valid_read ), 
	.D(n9522), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell4/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell4/controller/valid_read ), 
	.D(n9525), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell10/controller/valid_read ), 
	.D(n9531), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell4/reg_ptok/token_reg  (.RN(n3858), 
	.QN(\fifo_to_fft/hang[3] ), 
	.Q(n3994), 
	.D(n3993), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell4/reg_ptok/token_reg  (.RN(n4033), 
	.QN(\fifo_to_fir/hang[3] ), 
	.Q(n4169), 
	.D(n4168), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell2/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell2/reg_gtok/token ), 
	.D(n5508), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell2/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell2/reg_gtok/token ), 
	.D(n5560), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell8/reg_gtok/token ), 
	.D(n6752), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell8/reg_gtok/token ), 
	.D(n6223), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell3/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell3/controller/valid_read ), 
	.D(n9516), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell9/controller/valid_read ), 
	.D(n9522), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell3/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell3/controller/valid_read ), 
	.D(n9524), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell9/controller/valid_read ), 
	.D(n9529), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell9/reg_ptok/token_reg  (.RN(n4661), 
	.QN(\fifo_from_fir/hang[8] ), 
	.Q(n4802), 
	.D(n4801), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell2/reg_ptok/token_reg  (.RN(n3854), 
	.QN(\fifo_to_fft/hang[1] ), 
	.Q(n4000), 
	.D(n3999), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fft/fifo_cell3/reg_ptok/token_reg  (.RN(n3856), 
	.QN(\fifo_to_fft/hang[2] ), 
	.Q(n3997), 
	.D(n3996), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell2/reg_ptok/token_reg  (.RN(n4029), 
	.QN(\fifo_to_fir/hang[1] ), 
	.Q(n4175), 
	.D(n4174), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_to_fir/fifo_cell3/reg_ptok/token_reg  (.RN(n4031), 
	.QN(\fifo_to_fir/hang[2] ), 
	.Q(n4172), 
	.D(n4171), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell9/reg_ptok/token_reg  (.RN(n4475), 
	.QN(\fifo_from_fft/hang[8] ), 
	.Q(n4616), 
	.D(n4615), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/fir_put_req_reg  (.Q(\router/fir_put_req_reg ), 
	.D(n5459), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell1/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell1/reg_gtok/token ), 
	.D(n5511), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell1/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell1/reg_gtok/token ), 
	.D(n5563), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell1/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell1/controller/valid_read ), 
	.D(n9519), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell1/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell1/controller/valid_read ), 
	.D(n9524), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell1/reg_ptok/token_reg  (.Q(\fifo_to_fft/hang[0] ), 
	.D(n5517), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell1/reg_ptok/token_reg  (.Q(\fifo_to_fir/hang[0] ), 
	.D(n5569), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell2/controller/valid_read_reg  (.Q(\fifo_to_fft/fifo_cell2/controller/valid_read ), 
	.D(n9516), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell2/controller/valid_read_reg  (.Q(\fifo_to_fir/fifo_cell2/controller/valid_read ), 
	.D(n9524), 
	.CK(clk__L1_N0));
   EDFFTRX1TS \router/data_cntl/fft_put_req_reg  (.RN(n2848), 
	.QN(\router/fft_put_req_reg ), 
	.E(n3831), 
	.D(n7611), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell0/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell0/controller/f_i_get ), 
	.D(n5456), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell15/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell15/controller/f_i_get ), 
	.D(n5471), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell14/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell14/controller/f_i_get ), 
	.D(n5474), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell13/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell13/controller/f_i_get ), 
	.D(n5477), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell12/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell12/controller/f_i_get ), 
	.D(n5480), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell11/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell11/controller/f_i_get ), 
	.D(n5483), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell10/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell10/controller/f_i_get ), 
	.D(n5486), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell9/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell9/controller/f_i_get ), 
	.D(n5489), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell8/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell8/controller/f_i_get ), 
	.D(n5492), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell7/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell7/controller/f_i_get ), 
	.D(n5495), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell6/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell6/controller/f_i_get ), 
	.D(n5498), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell5/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell5/controller/f_i_get ), 
	.D(n5501), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell4/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell4/controller/f_i_get ), 
	.D(n5504), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell3/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell3/controller/f_i_get ), 
	.D(n5507), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell2/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell2/controller/f_i_get ), 
	.D(n5510), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell1/controller/f_i_get_reg  (.Q(\fifo_to_fft/fifo_cell1/controller/f_i_get ), 
	.D(n5513), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell0/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell0/controller/f_i_get ), 
	.D(n5454), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell1/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell1/controller/f_i_get ), 
	.D(n5565), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell0/reg_gtok/token_reg  (.Q(\fifo_to_fft/fifo_cell0/reg_gtok/token ), 
	.D(n5514), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell0/reg_gtok/token_reg  (.Q(\fifo_to_fir/fifo_cell0/reg_gtok/token ), 
	.D(n5566), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell7/reg_gtok/token ), 
	.D(n6753), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell7/reg_gtok/token ), 
	.D(n6224), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell0/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell0/controller/f_i_put ), 
	.D(n5515), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell14/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell14/controller/f_i_put ), 
	.D(n5473), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell13/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell13/controller/f_i_put ), 
	.D(n5476), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell12/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell12/controller/f_i_put ), 
	.D(n5479), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell10/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell10/controller/f_i_put ), 
	.D(n5485), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell9/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell9/controller/f_i_put ), 
	.D(n5488), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell8/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell8/controller/f_i_put ), 
	.D(n5491), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell6/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell6/controller/f_i_put ), 
	.D(n5497), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell5/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell5/controller/f_i_put ), 
	.D(n5500), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell4/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell4/controller/f_i_put ), 
	.D(n5503), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell3/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell3/controller/f_i_put ), 
	.D(n5506), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell2/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell2/controller/f_i_put ), 
	.D(n5509), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell1/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell1/controller/f_i_put ), 
	.D(n5512), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell8/controller/valid_read ), 
	.D(n9522), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell8/controller/valid_read ), 
	.D(n9530), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell8/reg_ptok/token_reg  (.RN(n4659), 
	.QN(\fifo_from_fir/hang[7] ), 
	.Q(n4805), 
	.D(n4804), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell8/reg_ptok/token_reg  (.RN(n4473), 
	.QN(\fifo_from_fft/hang[7] ), 
	.Q(n4619), 
	.D(n4618), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell15/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell15/controller/f_i_get ), 
	.D(n5523), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell14/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell14/controller/f_i_get ), 
	.D(n5526), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell13/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell13/controller/f_i_get ), 
	.D(n5529), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell12/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell12/controller/f_i_get ), 
	.D(n5532), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell11/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell11/controller/f_i_get ), 
	.D(n5535), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell10/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell10/controller/f_i_get ), 
	.D(n5538), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell9/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell9/controller/f_i_get ), 
	.D(n5541), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell8/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell8/controller/f_i_get ), 
	.D(n5544), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell7/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell7/controller/f_i_get ), 
	.D(n5547), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell6/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell6/controller/f_i_get ), 
	.D(n5550), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell5/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell5/controller/f_i_get ), 
	.D(n5553), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell4/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell4/controller/f_i_get ), 
	.D(n5556), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell3/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell3/controller/f_i_get ), 
	.D(n5559), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell2/controller/f_i_get_reg  (.Q(\fifo_to_fir/fifo_cell2/controller/f_i_get ), 
	.D(n5562), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell15/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell15/controller/f_i_put ), 
	.D(n5470), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell11/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell11/controller/f_i_put ), 
	.D(n5482), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fft/fifo_cell7/controller/f_i_put_reg  (.Q(\fifo_to_fft/fifo_cell7/controller/f_i_put ), 
	.D(n5494), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell0/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell0/controller/f_i_put ), 
	.D(n5567), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell15/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell15/controller/f_i_put ), 
	.D(n5522), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell14/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell14/controller/f_i_put ), 
	.D(n5525), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell13/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell13/controller/f_i_put ), 
	.D(n5528), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell12/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell12/controller/f_i_put ), 
	.D(n5531), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell11/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell11/controller/f_i_put ), 
	.D(n5534), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell10/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell10/controller/f_i_put ), 
	.D(n5537), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell9/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell9/controller/f_i_put ), 
	.D(n5540), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell8/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell8/controller/f_i_put ), 
	.D(n5543), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell7/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell7/controller/f_i_put ), 
	.D(n5546), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell6/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell6/controller/f_i_put ), 
	.D(n5549), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell5/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell5/controller/f_i_put ), 
	.D(n5552), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell4/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell4/controller/f_i_put ), 
	.D(n5555), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell3/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell3/controller/f_i_put ), 
	.D(n5558), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell2/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell2/controller/f_i_put ), 
	.D(n5561), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_to_fir/fifo_cell1/controller/f_i_put_reg  (.Q(\fifo_to_fir/fifo_cell1/controller/f_i_put ), 
	.D(n5564), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell7/controller/valid_read ), 
	.D(n9521), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell7/controller/valid_read ), 
	.D(n9530), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell7/reg_ptok/token_reg  (.RN(n4657), 
	.QN(\fifo_from_fir/hang[6] ), 
	.Q(n4808), 
	.D(n4807), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell7/reg_ptok/token_reg  (.RN(n4471), 
	.QN(\fifo_from_fft/hang[6] ), 
	.Q(n4622), 
	.D(n4621), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell6/reg_gtok/token ), 
	.D(n6754), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell6/reg_gtok/token ), 
	.D(n6225), 
	.CK(clk__L1_N0));
   DFFQX4TS \fifo_to_fft/empty_det/result_reg  (.Q(to_fft_empty), 
	.D(\fifo_to_fft/empty_det/N4 ), 
	.CK(clk__L1_N0));
   DFFQX4TS \fifo_to_fir/empty_det/result_reg  (.Q(to_fir_empty), 
	.D(\fifo_to_fir/empty_det/N4 ), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell6/reg_ptok/token_reg  (.RN(n4655), 
	.QN(\fifo_from_fir/hang[5] ), 
	.Q(n4811), 
	.D(n4810), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell6/reg_ptok/token_reg  (.RN(n4469), 
	.QN(\fifo_from_fft/hang[5] ), 
	.Q(n4625), 
	.D(n4624), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell5/reg_gtok/token ), 
	.D(n6755), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell5/reg_gtok/token ), 
	.D(n6226), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell6/controller/valid_read ), 
	.D(n9521), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell6/controller/valid_read ), 
	.D(n9529), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell4/reg_gtok/token ), 
	.D(n6756), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell4/reg_gtok/token ), 
	.D(n6227), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell5/controller/valid_read ), 
	.D(n9521), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell5/controller/valid_read ), 
	.D(n9530), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell5/reg_ptok/token_reg  (.RN(n4653), 
	.QN(\fifo_from_fir/hang[4] ), 
	.Q(n4814), 
	.D(n4813), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell5/reg_ptok/token_reg  (.RN(n4467), 
	.QN(\fifo_from_fft/hang[4] ), 
	.Q(n4628), 
	.D(n4627), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell3/reg_gtok/token ), 
	.D(n6757), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell3/reg_gtok/token ), 
	.D(n6228), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell4/controller/valid_read ), 
	.D(n9521), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell4/controller/valid_read ), 
	.D(n9530), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell4/reg_ptok/token_reg  (.RN(n4651), 
	.QN(\fifo_from_fir/hang[3] ), 
	.Q(n4817), 
	.D(n4816), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell4/reg_ptok/token_reg  (.RN(n4465), 
	.QN(\fifo_from_fft/hang[3] ), 
	.Q(n4631), 
	.D(n4630), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell3/controller/valid_read ), 
	.D(n9520), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell3/controller/valid_read ), 
	.D(n9528), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell3/reg_ptok/token_reg  (.RN(n4649), 
	.QN(\fifo_from_fir/hang[2] ), 
	.Q(n4820), 
	.D(n4819), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell3/reg_ptok/token_reg  (.RN(n4463), 
	.QN(\fifo_from_fft/hang[2] ), 
	.Q(n4634), 
	.D(n4633), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell2/reg_gtok/token ), 
	.D(n6758), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell2/reg_gtok/token ), 
	.D(n6229), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell2/reg_ptok/token_reg  (.RN(n4647), 
	.QN(\fifo_from_fir/hang[1] ), 
	.Q(n4823), 
	.D(n4822), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell1/reg_gtok/token ), 
	.D(n6759), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell1/reg_gtok/token ), 
	.D(n6230), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell2/controller/valid_read ), 
	.D(n9520), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell2/controller/valid_read ), 
	.D(n9528), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell2/reg_ptok/token_reg  (.RN(n4461), 
	.QN(\fifo_from_fft/hang[1] ), 
	.Q(n4637), 
	.D(n4636), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/reg_gtok/token_reg  (.Q(\fifo_from_fir/fifo_cell0/reg_gtok/token ), 
	.D(n6760), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/controller/valid_read_reg  (.Q(\fifo_from_fft/fifo_cell1/controller/valid_read ), 
	.D(n9520), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/controller/valid_read_reg  (.Q(\fifo_from_fir/fifo_cell1/controller/valid_read ), 
	.D(n9528), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fir/fifo_cell1/reg_ptok/token_reg  (.RN(n4645), 
	.QN(\fifo_from_fir/hang[0] ), 
	.Q(n4826), 
	.D(n4825), 
	.CK(clk__L1_N0));
   DFFTRX2TS \fifo_from_fft/fifo_cell1/reg_ptok/token_reg  (.RN(n4459), 
	.QN(\fifo_from_fft/hang[0] ), 
	.Q(n4640), 
	.D(n4639), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/fir_get_req_reg  (.Q(\router/fir_get_req_reg ), 
	.D(n6761), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/reg_gtok/token_reg  (.Q(\fifo_from_fft/fifo_cell0/reg_gtok/token ), 
	.D(n6231), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/pla_top/fir_enable_reg  (.Q(n9615), 
	.D(n5573), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/fir_read_calc/counter/done_reg  (.Q(\router/fir_read_done ), 
	.D(n5571), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/fir_write_calc/counter/done_reg  (.Q(\router/fir_write_done ), 
	.D(n5519), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/fft_write_calc/counter/done_reg  (.Q(\router/fft_write_done ), 
	.D(FE_OFN961_n5467), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/addr_calc/fft_read_calc/counter/done_reg  (.Q(\router/fft_read_done ), 
	.D(n5704), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/data_cntl/fft_get_req_reg  (.Q(\router/fft_get_req_reg ), 
	.D(n6232), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell0/controller/f_i_get ), 
	.D(n5417), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell1/controller/f_i_get ), 
	.D(n6742), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell2/controller/f_i_get ), 
	.D(n6708), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell3/controller/f_i_get ), 
	.D(n6674), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell4/controller/f_i_get ), 
	.D(n6640), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell5/controller/f_i_get ), 
	.D(n6606), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell6/controller/f_i_get ), 
	.D(n6572), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell7/controller/f_i_get ), 
	.D(n6538), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell8/controller/f_i_get ), 
	.D(n6504), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell9/controller/f_i_get ), 
	.D(n6470), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell10/controller/f_i_get ), 
	.D(n6436), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell11/controller/f_i_get ), 
	.D(n6402), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell12/controller/f_i_get ), 
	.D(n6368), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell13/controller/f_i_get ), 
	.D(n6334), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell14/controller/f_i_get ), 
	.D(n6300), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/controller/f_i_get_reg  (.Q(\fifo_from_fir/fifo_cell15/controller/f_i_get ), 
	.D(n6266), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/pla_top/fft_enable_reg  (.Q(n9614), 
	.D(n5466), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell0/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell0/controller/f_i_put ), 
	.D(n6744), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell1/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell1/controller/f_i_put ), 
	.D(n6743), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell2/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell2/controller/f_i_put ), 
	.D(n6709), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell3/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell3/controller/f_i_put ), 
	.D(n6675), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell4/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell4/controller/f_i_put ), 
	.D(n6641), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell5/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell5/controller/f_i_put ), 
	.D(n6607), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell6/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell6/controller/f_i_put ), 
	.D(n6573), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell7/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell7/controller/f_i_put ), 
	.D(n6539), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell8/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell8/controller/f_i_put ), 
	.D(n6505), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell9/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell9/controller/f_i_put ), 
	.D(n6471), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell10/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell10/controller/f_i_put ), 
	.D(n6437), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell11/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell11/controller/f_i_put ), 
	.D(n6403), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell12/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell12/controller/f_i_put ), 
	.D(n6369), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell13/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell13/controller/f_i_put ), 
	.D(n6335), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell14/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell14/controller/f_i_put ), 
	.D(n6301), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fir/fifo_cell15/controller/f_i_put_reg  (.Q(\fifo_from_fir/fifo_cell15/controller/f_i_put ), 
	.D(n6267), 
	.CK(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[31]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[31] ), 
	.D(n5574), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[30]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[30] ), 
	.D(n5575), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[29]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[29] ), 
	.D(n5576), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[28]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[28] ), 
	.D(n5577), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[27]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[27] ), 
	.D(n5578), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[26]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[26] ), 
	.D(n5579), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[0]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[0] ), 
	.D(n5605), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[1]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[1] ), 
	.D(n5604), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[2]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[2] ), 
	.D(n5603), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[3]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[3] ), 
	.D(n5602), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[4]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[4] ), 
	.D(n5601), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[5]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[5] ), 
	.D(n5600), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[6]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[6] ), 
	.D(n5599), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[7]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[7] ), 
	.D(n5598), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[8]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[8] ), 
	.D(n5597), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[9]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[9] ), 
	.D(n5596), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[10]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[10] ), 
	.D(n5595), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[11]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[11] ), 
	.D(n5594), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[12]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[12] ), 
	.D(n5593), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[13]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[13] ), 
	.D(n5592), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[14]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[14] ), 
	.D(n5591), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[15]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[15] ), 
	.D(n5590), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[16]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[16] ), 
	.D(n5589), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[17]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[17] ), 
	.D(n5588), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[18]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[18] ), 
	.D(n5587), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[19]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[19] ), 
	.D(n5586), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[20]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[20] ), 
	.D(n5585), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[21]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[21] ), 
	.D(n5584), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[22]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[22] ), 
	.D(n5583), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[23]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[23] ), 
	.D(n5582), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[24]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[24] ), 
	.D(n5581), 
	.CKN(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accfullinstruction_reg[25]  (.SN(1'b1), 
	.RN(1'b1), 
	.Q(\mips/mips/accfullinstruction[25] ), 
	.D(n5580), 
	.CKN(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell0/controller/f_i_get ), 
	.D(n5452), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell1/controller/f_i_get ), 
	.D(n6213), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell2/controller/f_i_get ), 
	.D(n6179), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell3/controller/f_i_get ), 
	.D(n6145), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell4/controller/f_i_get ), 
	.D(n6111), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell5/controller/f_i_get ), 
	.D(n6077), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell6/controller/f_i_get ), 
	.D(n6043), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell7/controller/f_i_get ), 
	.D(n6009), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell8/controller/f_i_get ), 
	.D(n5975), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell9/controller/f_i_get ), 
	.D(n5941), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell10/controller/f_i_get ), 
	.D(n5907), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell11/controller/f_i_get ), 
	.D(n5873), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell12/controller/f_i_get ), 
	.D(n5839), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell13/controller/f_i_get ), 
	.D(n5805), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell14/controller/f_i_get ), 
	.D(n5771), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/controller/f_i_get_reg  (.Q(\fifo_from_fft/fifo_cell15/controller/f_i_get ), 
	.D(n5737), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell0/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell0/controller/f_i_put ), 
	.D(n6215), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell1/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell1/controller/f_i_put ), 
	.D(n6214), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell2/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell2/controller/f_i_put ), 
	.D(n6180), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell3/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell3/controller/f_i_put ), 
	.D(n6146), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell4/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell4/controller/f_i_put ), 
	.D(n6112), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell5/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell5/controller/f_i_put ), 
	.D(n6078), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell6/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell6/controller/f_i_put ), 
	.D(n6044), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell7/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell7/controller/f_i_put ), 
	.D(n6010), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell8/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell8/controller/f_i_put ), 
	.D(n5976), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell9/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell9/controller/f_i_put ), 
	.D(n5942), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell10/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell10/controller/f_i_put ), 
	.D(n5908), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell11/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell11/controller/f_i_put ), 
	.D(n5874), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell12/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell12/controller/f_i_put ), 
	.D(n5840), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell13/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell13/controller/f_i_put ), 
	.D(n5806), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell14/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell14/controller/f_i_put ), 
	.D(n5772), 
	.CK(clk__L1_N0));
   DFFQX1TS \fifo_from_fft/fifo_cell15/controller/f_i_put_reg  (.Q(\fifo_from_fft/fifo_cell15/controller/f_i_put ), 
	.D(n5738), 
	.CK(clk__L1_N0));
   DFFQX1TS \router/pla_top/acc_done_reg  (.Q(acc_done), 
	.D(n5703), 
	.CK(clk__L1_N0));
   DFFNSRX2TS \mips/mips/c/md/accbypass_reg  (.SN(1'b1), 
	.RN(1'b1), 
	.QN(n4311), 
	.Q(\mips/mips/accbypass ), 
	.D(n5702), 
	.CKN(clk__L1_N0));
   INVX2TS U3842 (.Y(\fifo_from_fft/fifo_cell15/data_out/N35 ), 
	.A(n4494));
   INVX2TS U3836 (.Y(\fifo_from_fft/fifo_cell14/data_out/N35 ), 
	.A(n4500));
   INVX2TS U3854 (.Y(\fifo_from_fft/fifo_cell13/data_out/N35 ), 
	.A(n4506));
   INVX2TS U3856 (.Y(\fifo_from_fft/fifo_cell1/data_out/N35 ), 
	.A(n4578));
   INVX2TS U3699 (.Y(\fifo_from_fir/fifo_cell15/data_out/N35 ), 
	.A(n4680));
   INVX2TS U3693 (.Y(\fifo_from_fir/fifo_cell14/data_out/N35 ), 
	.A(n4686));
   INVX2TS U3711 (.Y(\fifo_from_fir/fifo_cell13/data_out/N35 ), 
	.A(n4692));
   INVX2TS U3713 (.Y(\fifo_from_fir/fifo_cell1/data_out/N35 ), 
	.A(n4764));
   OAI21XLTS U1421 (.Y(n4443), 
	.B0(n4444), 
	.A1(n4442), 
	.A0(n4441));
   INVX2TS U3383 (.Y(\fifo_to_fir/fifo_cell2/data_out/N35 ), 
	.A(n4123));
   INVX2TS U3412 (.Y(\fifo_to_fir/fifo_cell4/data_out/N35 ), 
	.A(n4113));
   INVX2TS U3526 (.Y(\fifo_to_fft/fifo_cell2/data_out/N35 ), 
	.A(n3948));
   AOI22XLTS U347 (.Y(n3551), 
	.B1(\router/addr_calc/fir_write_calc/counter/N57 ), 
	.B0(FE_OFN892_n3531), 
	.A1(FE_OFN907_n3530), 
	.A0(n7205));
   AOI22XLTS U351 (.Y(n3553), 
	.B1(\router/addr_calc/fir_write_calc/counter/N55 ), 
	.B0(FE_OFN889_n3531), 
	.A1(FE_OFN904_n3530), 
	.A0(FE_OFN1266_router_addr_calc_fir_write_calc_count_9_));
   AOI22XLTS U576 (.Y(n3685), 
	.B1(\router/addr_calc/fft_read_calc/counter/N55 ), 
	.B0(FE_OFN867_n3663), 
	.A1(FE_OFN885_n3662), 
	.A0(FE_OFN1267_router_addr_calc_fft_read_calc_count_9_));
   AOI22XLTS U572 (.Y(n3683), 
	.B1(\router/addr_calc/fft_read_calc/counter/N57 ), 
	.B0(FE_OFN869_n3663), 
	.A1(FE_OFN885_n3662), 
	.A0(n7561));
   AOI22XLTS U426 (.Y(n3597), 
	.B1(\router/addr_calc/fir_read_calc/counter/N55 ), 
	.B0(n3575), 
	.A1(FE_OFN921_n3574), 
	.A0(\router/addr_calc/fir_read_calc/count[9] ));
   AOI22XLTS U501 (.Y(n3641), 
	.B1(\router/addr_calc/fft_write_calc/counter/N55 ), 
	.B0(FE_OFN958_n3619), 
	.A1(FE_OFN965_n3618), 
	.A0(FE_OFN1268_router_addr_calc_fft_write_calc_count_9_));
   AOI22XLTS U422 (.Y(n3595), 
	.B1(\router/addr_calc/fir_read_calc/counter/N57 ), 
	.B0(FE_OFN912_n3575), 
	.A1(FE_OFN923_n3574), 
	.A0(n7323));
   AOI22XLTS U497 (.Y(n3639), 
	.B1(\router/addr_calc/fft_write_calc/counter/N57 ), 
	.B0(FE_OFN957_n3619), 
	.A1(FE_OFN965_n3618), 
	.A0(n7437));
   AOI22XLTS U475 (.Y(n3628), 
	.B1(\router/addr_calc/fft_write_calc/counter/N68 ), 
	.B0(FE_OFN955_n3619), 
	.A1(FE_OFN969_n3618), 
	.A0(FE_OFN1249_n7392));
   AOI22XLTS U400 (.Y(n3584), 
	.B1(\router/addr_calc/fir_read_calc/counter/N68 ), 
	.B0(FE_OFN916_n3575), 
	.A1(FE_OFN927_n3574), 
	.A0(FE_OFN1250_n7278));
   AOI22XLTS U325 (.Y(n3540), 
	.B1(\router/addr_calc/fir_write_calc/counter/N68 ), 
	.B0(FE_OFN891_n3531), 
	.A1(FE_OFN905_n3530), 
	.A0(FE_OFN1251_n7153));
   AOI22XLTS U550 (.Y(n3672), 
	.B1(\router/addr_calc/fft_read_calc/counter/N68 ), 
	.B0(FE_OFN874_n3663), 
	.A1(FE_OFN883_n3662), 
	.A0(n7516));
   AOI22XLTS U329 (.Y(n3542), 
	.B1(\router/addr_calc/fir_write_calc/counter/N66 ), 
	.B0(FE_OFN895_n3531), 
	.A1(FE_OFN905_n3530), 
	.A0(FE_OFN1257_n7165));
   AOI22XLTS U554 (.Y(n3674), 
	.B1(\router/addr_calc/fft_read_calc/counter/N66 ), 
	.B0(FE_OFN874_n3663), 
	.A1(FE_OFN884_n3662), 
	.A0(n7526));
   AOI22XLTS U479 (.Y(n3630), 
	.B1(\router/addr_calc/fft_write_calc/counter/N66 ), 
	.B0(FE_OFN953_n3619), 
	.A1(FE_OFN968_n3618), 
	.A0(FE_OFN1255_n7402));
   AOI22XLTS U404 (.Y(n3586), 
	.B1(\router/addr_calc/fir_read_calc/counter/N66 ), 
	.B0(FE_OFN915_n3575), 
	.A1(FE_OFN926_n3574), 
	.A0(FE_OFN1256_n7288));
   AOI22XLTS U278 (.Y(n3510), 
	.B1(\router/addr_calc/iir_write_calc/counter/N54 ), 
	.B0(FE_OFN936_n3487), 
	.A1(FE_OFN947_n3486), 
	.A0(n7098));
   AOI22XLTS U288 (.Y(n3515), 
	.B1(\router/addr_calc/iir_write_calc/counter/N49 ), 
	.B0(FE_OFN939_n3487), 
	.A1(FE_OFN942_n3486), 
	.A0(n7101));
   AOI22XLTS U272 (.Y(n3507), 
	.B1(\router/addr_calc/iir_write_calc/counter/N57 ), 
	.B0(FE_OFN935_n3487), 
	.A1(FE_OFN948_n3486), 
	.A0(n7109));
   NOR3XLTS U957 (.Y(n5520), 
	.C(FE_OFN991_n9431), 
	.B(n3530), 
	.A(\router/addr_calc/fir_write_calc/counter/hold ));
   NOR3XLTS U784 (.Y(n5457), 
	.C(FE_OFN974_n9462), 
	.B(FE_OFN878_n3662), 
	.A(\router/addr_calc/fft_read_calc/counter/hold ));
   NOR3XLTS U813 (.Y(n5468), 
	.C(FE_OFN982_n9462), 
	.B(n3618), 
	.A(\router/addr_calc/fft_write_calc/counter/hold ));
   NOR3XLTS U1101 (.Y(n5572), 
	.C(n9431), 
	.B(FE_OFN929_n3574), 
	.A(\router/addr_calc/fir_read_calc/counter/hold ));
   NOR3XLTS U612 (.Y(n3712), 
	.C(n3716), 
	.B(n9434), 
	.A(FE_OFN1283_router_fft_write_done));
   AOI211XLTS U609 (.Y(n3709), 
	.C0(n3710), 
	.B0(n9389), 
	.A1(\router/fir_write_done ), 
	.A0(n9406));
   OAI32XLTS U1099 (.Y(n5571), 
	.B1(FE_OFN1190_n7022), 
	.B0(n7211), 
	.A2(FE_OFN985_n9431), 
	.A1(\router/addr_calc/fir_read_calc/counter/N40 ), 
	.A0(\router/addr_calc/fir_read_calc/counter/hold ));
   OAI32X1TS U811 (.Y(n5467), 
	.B1(n7019), 
	.B0(n3850), 
	.A2(FE_OFN981_n9462), 
	.A1(\router/addr_calc/fft_write_calc/counter/N40 ), 
	.A0(\router/addr_calc/fft_write_calc/counter/hold ));
   INVXLTS U1442 (.Y(n4458), 
	.A(\router/fft_read_done ));
   OAI32X1TS U1440 (.Y(n5704), 
	.B1(FE_OFN1168_n7021), 
	.B0(n4458), 
	.A2(n9462), 
	.A1(\router/addr_calc/fft_read_calc/counter/N40 ), 
	.A0(\router/addr_calc/fft_read_calc/counter/hold ));
   OAI32X1TS U955 (.Y(n5519), 
	.B1(n7020), 
	.B0(n4025), 
	.A2(FE_OFN991_n9431), 
	.A1(\router/addr_calc/fir_write_calc/counter/N40 ), 
	.A0(\router/addr_calc/fir_write_calc/counter/hold ));
   AOI21XLTS U788 (.Y(n3824), 
	.B0(n3825), 
	.A1(\router/fir_put_req_reg ), 
	.A0(n3823));
   NOR3XLTS U2752 (.Y(n6766), 
	.C(n9389), 
	.B(n3486), 
	.A(\router/addr_calc/iir_write_calc/counter/hold ));
   OAI21XLTS U1436 (.Y(n3849), 
	.B0(n4455), 
	.A1(n3850), 
	.A0(n7960));
   OAI211XLTS U1435 (.Y(n4450), 
	.C0(n3849), 
	.B0(acc_done), 
	.A1(n4457), 
	.A0(n4203));
   AND3XLTS U3616 (.Y(\fifo_from_fir/fifo_cell15/N7 ), 
	.C(\fifo_from_fir/fifo_cell15/data_out/N9 ), 
	.B(FE_OFN742_n4829), 
	.A(\fifo_from_fir/fifo_cell15/reg_gtok/token ));
   OAI32X1TS U2749 (.Y(n6765), 
	.B1(\router/addr_calc/iir_write_calc/counter/N212 ), 
	.B0(n3717), 
	.A2(n9389), 
	.A1(\router/addr_calc/iir_write_calc/counter/N40 ), 
	.A0(\router/addr_calc/iir_write_calc/counter/hold ));
   OAI31X1TS U809 (.Y(n5466), 
	.B0(n3847), 
	.A2(n3846), 
	.A1(FE_OFN1283_router_fft_write_done), 
	.A0(FE_OFN839_n7619));
   AND2XLTS U801 (.Y(n5461), 
	.B(n3839), 
	.A(\router/data_cntl/N151 ));
   AOI31XLTS U793 (.Y(n3833), 
	.B0(n3830), 
	.A2(FE_OFN1284_router_ram_read_enable_reg), 
	.A1(n9434), 
	.A0(n3476));
   MX2XLTS U792 (.Y(n5460), 
	.S0(n3833), 
	.B(\router/data_cntl/fft_full_flag ), 
	.A(FE_OFN1284_router_ram_read_enable_reg));
   OAI32XLTS U804 (.Y(n5464), 
	.B1(n3844), 
	.B0(\router/addr_calc/N95 ), 
	.A2(n3843), 
	.A1(n7207), 
	.A0(n3842));
   AND3XLTS U3759 (.Y(\fifo_from_fft/fifo_cell15/N7 ), 
	.C(\fifo_from_fft/fifo_cell15/data_out/N9 ), 
	.B(FE_OFN724_n4643), 
	.A(\fifo_from_fft/fifo_cell15/reg_gtok/token ));
   OAI22XLTS U806 (.Y(n5465), 
	.B1(n3844), 
	.B0(\router/addr_calc/N99 ), 
	.A1(n7207), 
	.A0(n3845));
   AOI211XLTS U803 (.Y(n5463), 
	.C0(n3841), 
	.B0(FE_OFN981_n9462), 
	.A1(\router/addr_calc/N9 ), 
	.A0(FE_OFN1438_router_data_from_fft));
   AOI211XLTS U802 (.Y(n5462), 
	.C0(n3840), 
	.B0(FE_OFN980_n9462), 
	.A1(\router/addr_calc/N63 ), 
	.A0(\router/data_to_fft ));
   OAI32XLTS U216 (.Y(\router/data_cntl/N139 ), 
	.B1(n3463), 
	.B0(to_fir_empty), 
	.A2(n3465), 
	.A1(n3474), 
	.A0(n3463));
   OAI211X1TS U215 (.Y(\router/data_cntl/N142 ), 
	.C0(FE_OFN990_n9431), 
	.B0(FE_OFN977_n9462), 
	.A1(n9390), 
	.A0(FE_OFN1285_router_ram_read_enable_reg));
   OAI21XLTS U3317 (.Y(\mips/mips/a/N50 ), 
	.B0(n4444), 
	.A1(n4445), 
	.A0(n4441));
   INVX2TS U3321 (.Y(\mips/mips/a/N49 ), 
	.A(n4444));
   INVX2TS U1427 (.Y(n3456), 
	.A(n4205));
   INVX2TS U3813 (.Y(n4641), 
	.A(n4460));
   INVX2TS U3804 (.Y(n4635), 
	.A(n4464));
   INVX2TS U3800 (.Y(n4632), 
	.A(n4466));
   INVX2TS U3796 (.Y(n4629), 
	.A(n4468));
   INVX2TS U3792 (.Y(n4626), 
	.A(n4470));
   INVX2TS U3788 (.Y(n4623), 
	.A(n4472));
   INVX2TS U3784 (.Y(n4620), 
	.A(n4474));
   INVX2TS U3780 (.Y(n4617), 
	.A(n4476));
   INVX2TS U3776 (.Y(n4614), 
	.A(n4478));
   INVX2TS U3772 (.Y(n4611), 
	.A(n4480));
   INVX2TS U3768 (.Y(n4608), 
	.A(n4482));
   INVX2TS U3764 (.Y(n4605), 
	.A(n4484));
   INVX2TS U3760 (.Y(n4602), 
	.A(n4486));
   NOR2X1TS U735 (.Y(n3788), 
	.B(n8845), 
	.A(n3787));
   OAI32X1TS U732 (.Y(n5419), 
	.B1(n3791), 
	.B0(n8840), 
	.A2(n3789), 
	.A1(FE_OFN783_n7619), 
	.A0(n3788));
   INVX2TS U3670 (.Y(n4827), 
	.A(n4646));
   INVX2TS U3661 (.Y(n4821), 
	.A(n4650));
   INVX2TS U3657 (.Y(n4818), 
	.A(n4652));
   INVX2TS U3653 (.Y(n4815), 
	.A(n4654));
   INVX2TS U3649 (.Y(n4812), 
	.A(n4656));
   INVX2TS U3645 (.Y(n4809), 
	.A(n4658));
   INVX2TS U3641 (.Y(n4806), 
	.A(n4660));
   INVX2TS U3637 (.Y(n4803), 
	.A(n4662));
   INVX2TS U3633 (.Y(n4800), 
	.A(n4664));
   INVX2TS U3629 (.Y(n4797), 
	.A(n4666));
   INVX2TS U3625 (.Y(n4794), 
	.A(n4668));
   INVX2TS U3621 (.Y(n4791), 
	.A(n4670));
   INVX2TS U3617 (.Y(n4788), 
	.A(n4672));
   NOR2X1TS U689 (.Y(n3768), 
	.B(n8878), 
	.A(n3767));
   OAI32X1TS U686 (.Y(n5384), 
	.B1(n3771), 
	.B0(n8873), 
	.A2(n3769), 
	.A1(FE_OFN804_n7619), 
	.A0(n3768));
   OAI21X1TS U2000 (.Y(n3798), 
	.B0(n3796), 
	.A1(n4580), 
	.A0(n7222));
   AOI21X1TS U773 (.Y(n5452), 
	.B0(n7619), 
	.A1(n3798), 
	.A0(\fifo_from_fft/fifo_cell0/controller/valid_read ));
   OAI21X1TS U1999 (.Y(n6215), 
	.B0(n3798), 
	.A1(\fifo_from_fft/fifo_cell0/data_out/N35 ), 
	.A0(n4579));
   OAI21X1TS U2631 (.Y(n3778), 
	.B0(n3776), 
	.A1(n4766), 
	.A0(n7217));
   AOI21X1TS U727 (.Y(n5417), 
	.B0(FE_OFN809_n7619), 
	.A1(n3778), 
	.A0(\fifo_from_fir/fifo_cell0/controller/valid_read ));
   OAI21X1TS U2630 (.Y(n6744), 
	.B0(n3778), 
	.A1(\fifo_from_fir/fifo_cell0/data_out/N35 ), 
	.A0(n4765));
   OAI211X1TS U2024 (.Y(n4597), 
	.C0(n9473), 
	.B0(\fifo_from_fft/hang[14] ), 
	.A1(n4599), 
	.A0(n8840));
   AOI21X1TS U1477 (.Y(n5737), 
	.B0(FE_OFN802_n7619), 
	.A1(n4491), 
	.A0(\fifo_from_fft/fifo_cell15/controller/valid_read ));
   OAI211X1TS U2655 (.Y(n4783), 
	.C0(n9469), 
	.B0(\fifo_from_fir/hang[14] ), 
	.A1(n4785), 
	.A0(n8873));
   AOI21X1TS U1514 (.Y(n5771), 
	.B0(FE_OFN802_n7619), 
	.A1(n4497), 
	.A0(\fifo_from_fft/fifo_cell14/controller/valid_read ));
   AOI21X1TS U2108 (.Y(n6266), 
	.B0(FE_OFN788_n7619), 
	.A1(n4677), 
	.A0(\fifo_from_fir/fifo_cell15/controller/valid_read ));
   AOI21X1TS U2145 (.Y(n6300), 
	.B0(FE_OFN785_n7619), 
	.A1(n4683), 
	.A0(\fifo_from_fir/fifo_cell14/controller/valid_read ));
   AOI21X1TS U1551 (.Y(n5805), 
	.B0(FE_OFN802_n7619), 
	.A1(n4503), 
	.A0(\fifo_from_fft/fifo_cell13/controller/valid_read ));
   AOI21X1TS U2182 (.Y(n6334), 
	.B0(FE_OFN788_n7619), 
	.A1(n4689), 
	.A0(\fifo_from_fir/fifo_cell13/controller/valid_read ));
   AOI21X1TS U1588 (.Y(n5839), 
	.B0(FE_OFN806_n7619), 
	.A1(n4509), 
	.A0(\fifo_from_fft/fifo_cell12/controller/valid_read ));
   AOI21X1TS U2219 (.Y(n6368), 
	.B0(FE_OFN815_n7619), 
	.A1(n4695), 
	.A0(\fifo_from_fir/fifo_cell12/controller/valid_read ));
   INVX2TS U3368 (.Y(n4167), 
	.A(n4036));
   INVX2TS U3356 (.Y(n4158), 
	.A(n4042));
   INVX2TS U3344 (.Y(n4149), 
	.A(n4048));
   INVX2TS U3340 (.Y(n4146), 
	.A(n4050));
   INVX2TS U3398 (.Y(\fifo_to_fir/fifo_cell0/data_out/N35 ), 
	.A(n4133));
   OAI31X1TS U1075 (.Y(n3807), 
	.B0(\fifo_to_fir/fifo_cell0/reg_ptok/N29 ), 
	.A2(\fifo_to_fir/fifo_cell0/reg_ptok/N22 ), 
	.A1(\fifo_to_fir/fifo_cell0/reg_ptok/out_valid_get ), 
	.A0(\fifo_to_fir/fifo_cell0/reg_ptok/out_valid_put ));
   NOR3X1TS U3517 (.Y(n5244), 
	.C(\fifo_to_fft/fifo_cell4/controller/valid_read ), 
	.B(\fifo_to_fft/fifo_cell4/controller/write_enable ), 
	.A(n7321));
   INVX2TS U3511 (.Y(n3992), 
	.A(n3861));
   INVX2TS U3499 (.Y(n3983), 
	.A(n3867));
   INVX2TS U3487 (.Y(n3974), 
	.A(n3873));
   INVX2TS U3483 (.Y(n3971), 
	.A(n3875));
   INVX2TS U3479 (.Y(n3968), 
	.A(n3877));
   INVX2TS U3542 (.Y(\fifo_to_fft/fifo_cell0/data_out/N35 ), 
	.A(n3958));
   OAI31X1TS U931 (.Y(n3818), 
	.B0(\fifo_to_fft/fifo_cell0/reg_ptok/N29 ), 
	.A2(\fifo_to_fft/fifo_cell0/reg_ptok/N22 ), 
	.A1(\fifo_to_fft/fifo_cell0/reg_ptok/out_valid_get ), 
	.A0(\fifo_to_fft/fifo_cell0/reg_ptok/out_valid_put ));
   NOR2X1TS U930 (.Y(n4003), 
	.B(n8812), 
	.A(n3818));
   OAI21X1TS U928 (.Y(n4005), 
	.B0(n9496), 
	.A1(n3815), 
	.A0(n3814));
   OAI32X1TS U927 (.Y(n5518), 
	.B1(n4005), 
	.B0(n8808), 
	.A2(n4004), 
	.A1(FE_OFN786_n7619), 
	.A0(n4003));
   NOR2X1TS U1074 (.Y(n4178), 
	.B(n8791), 
	.A(n3807));
   OAI21X1TS U1072 (.Y(n4180), 
	.B0(n9496), 
	.A1(n3804), 
	.A0(n3803));
   OAI32X1TS U1071 (.Y(n5570), 
	.B1(n4180), 
	.B0(n8787), 
	.A2(n4179), 
	.A1(FE_OFN787_n7619), 
	.A0(n4178));
   AOI21X1TS U1033 (.Y(n5565), 
	.B0(FE_OFN779_n7619), 
	.A1(n4130), 
	.A0(\fifo_to_fir/fifo_cell1/controller/valid_read ));
   AOI21X1TS U889 (.Y(n5513), 
	.B0(FE_OFN794_n7619), 
	.A1(n3955), 
	.A0(\fifo_to_fft/fifo_cell1/controller/valid_read ));
   OAI21X1TS U887 (.Y(n5512), 
	.B0(n3955), 
	.A1(n3954), 
	.A0(\fifo_to_fft/fifo_cell1/data_out/N35 ));
   OAI21X1TS U1031 (.Y(n5564), 
	.B0(n4130), 
	.A1(n4129), 
	.A0(\fifo_to_fir/fifo_cell1/data_out/N35 ));
   OAI21X1TS U1038 (.Y(n3808), 
	.B0(n4136), 
	.A1(n4133), 
	.A0(n7227));
   OAI21X1TS U894 (.Y(n3819), 
	.B0(n3961), 
	.A1(n3958), 
	.A0(n7232));
   AOI21X1TS U783 (.Y(n5456), 
	.B0(FE_OFN782_n7619), 
	.A1(n3819), 
	.A0(\fifo_to_fft/fifo_cell0/controller/valid_read ));
   OAI21X1TS U1037 (.Y(n5567), 
	.B0(n3808), 
	.A1(\fifo_to_fir/fifo_cell0/data_out/N35 ), 
	.A0(n4135));
   OAI21X1TS U893 (.Y(n5515), 
	.B0(n3819), 
	.A1(\fifo_to_fft/fifo_cell0/data_out/N35 ), 
	.A0(n3960));
   OAI211X1TS U1041 (.Y(n4137), 
	.C0(n9476), 
	.B0(\fifo_to_fir/hang[14] ), 
	.A1(n4055), 
	.A0(n8789));
   OAI21X1TS U964 (.Y(n4060), 
	.B0(n4062), 
	.A1(n7346), 
	.A0(n7351));
   AOI21X1TS U963 (.Y(n5523), 
	.B0(FE_OFN798_n7619), 
	.A1(n4060), 
	.A0(\fifo_to_fir/fifo_cell15/controller/valid_read ));
   OAI21X1TS U820 (.Y(n3885), 
	.B0(n3887), 
	.A1(n7237), 
	.A0(n7242));
   AOI21X1TS U819 (.Y(n5471), 
	.B0(FE_OFN792_n7619), 
	.A1(n3885), 
	.A0(\fifo_to_fft/fifo_cell15/controller/valid_read ));
   OAI21X1TS U817 (.Y(n5470), 
	.B0(n3885), 
	.A1(n3884), 
	.A0(\fifo_to_fft/fifo_cell15/data_out/N35 ));
   OAI21X1TS U961 (.Y(n5522), 
	.B0(n4060), 
	.A1(n4059), 
	.A0(\fifo_to_fir/fifo_cell15/data_out/N35 ));
   AOI21X1TS U824 (.Y(n5474), 
	.B0(FE_OFN796_n7619), 
	.A1(n3890), 
	.A0(\fifo_to_fft/fifo_cell14/controller/valid_read ));
   AOI21X1TS U968 (.Y(n5526), 
	.B0(FE_OFN805_n7619), 
	.A1(n4065), 
	.A0(\fifo_to_fir/fifo_cell14/controller/valid_read ));
   OAI21X1TS U822 (.Y(n5473), 
	.B0(n3890), 
	.A1(n3889), 
	.A0(\fifo_to_fft/fifo_cell14/data_out/N35 ));
   OAI21X1TS U966 (.Y(n5525), 
	.B0(n4065), 
	.A1(n4064), 
	.A0(\fifo_to_fir/fifo_cell14/data_out/N35 ));
   OAI21X1TS U974 (.Y(n4070), 
	.B0(n7366), 
	.A1(n4068), 
	.A0(n7361));
   AOI21X1TS U973 (.Y(n5529), 
	.B0(FE_OFN814_n7619), 
	.A1(n4070), 
	.A0(\fifo_to_fir/fifo_cell13/controller/valid_read ));
   OAI21X1TS U830 (.Y(n3895), 
	.B0(n7256), 
	.A1(n3893), 
	.A0(n7252));
   AOI21X1TS U829 (.Y(n5477), 
	.B0(FE_OFN801_n7619), 
	.A1(n3895), 
	.A0(\fifo_to_fft/fifo_cell13/controller/valid_read ));
   OAI21X1TS U971 (.Y(n5528), 
	.B0(n4070), 
	.A1(n4069), 
	.A0(\fifo_to_fir/fifo_cell13/data_out/N35 ));
   OAI21X1TS U827 (.Y(n5476), 
	.B0(n3895), 
	.A1(n3894), 
	.A0(\fifo_to_fft/fifo_cell13/data_out/N35 ));
   OAI21X1TS U979 (.Y(n4075), 
	.B0(n7375), 
	.A1(n4073), 
	.A0(n7370));
   AOI21X1TS U978 (.Y(n5532), 
	.B0(FE_OFN810_n7619), 
	.A1(n4075), 
	.A0(\fifo_to_fir/fifo_cell12/controller/valid_read ));
   OAI21X1TS U835 (.Y(n3900), 
	.B0(n7266), 
	.A1(n3898), 
	.A0(n7261));
   AOI21X1TS U834 (.Y(n5480), 
	.B0(FE_OFN813_n7619), 
	.A1(n3900), 
	.A0(\fifo_to_fft/fifo_cell12/controller/valid_read ));
   OAI21X1TS U976 (.Y(n5531), 
	.B0(n4075), 
	.A1(n4074), 
	.A0(\fifo_to_fir/fifo_cell12/data_out/N35 ));
   OAI21X1TS U832 (.Y(n5479), 
	.B0(n3900), 
	.A1(n3899), 
	.A0(\fifo_to_fft/fifo_cell12/data_out/N35 ));
   AOI21X1TS U839 (.Y(n5483), 
	.B0(FE_OFN842_n7619), 
	.A1(n3905), 
	.A0(\fifo_to_fft/fifo_cell11/controller/valid_read ));
   AOI21X1TS U983 (.Y(n5535), 
	.B0(FE_OFN816_n7619), 
	.A1(n4080), 
	.A0(\fifo_to_fir/fifo_cell11/controller/valid_read ));
   OAI21X1TS U837 (.Y(n5482), 
	.B0(n3905), 
	.A1(n3904), 
	.A0(\fifo_to_fft/fifo_cell11/data_out/N35 ));
   OAI21X1TS U981 (.Y(n5534), 
	.B0(n4080), 
	.A1(n4079), 
	.A0(\fifo_to_fir/fifo_cell11/data_out/N35 ));
   OAI21X1TS U994 (.Y(n4090), 
	.B0(n7395), 
	.A1(n4088), 
	.A0(n7390));
   AOI21X1TS U993 (.Y(n5541), 
	.B0(FE_OFN823_n7619), 
	.A1(n4090), 
	.A0(\fifo_to_fir/fifo_cell9/controller/valid_read ));
   OAI21X1TS U850 (.Y(n3915), 
	.B0(n7286), 
	.A1(n3913), 
	.A0(n7281));
   AOI21X1TS U849 (.Y(n5489), 
	.B0(FE_OFN838_n7619), 
	.A1(n3915), 
	.A0(\fifo_to_fft/fifo_cell9/controller/valid_read ));
   OAI21X1TS U999 (.Y(n4095), 
	.B0(n7405), 
	.A1(n4093), 
	.A0(n7400));
   AOI21X1TS U998 (.Y(n5544), 
	.B0(FE_OFN823_n7619), 
	.A1(n4095), 
	.A0(\fifo_to_fir/fifo_cell8/controller/valid_read ));
   OAI21X1TS U855 (.Y(n3920), 
	.B0(FE_OFN678_n7295), 
	.A1(n3918), 
	.A0(n7291));
   AOI21X1TS U854 (.Y(n5492), 
	.B0(FE_OFN838_n7619), 
	.A1(n3920), 
	.A0(\fifo_to_fft/fifo_cell8/controller/valid_read ));
   OAI21X1TS U1009 (.Y(n4105), 
	.B0(n4107), 
	.A1(n4103), 
	.A0(n7415));
   OAI21X1TS U865 (.Y(n3930), 
	.B0(n3932), 
	.A1(n3928), 
	.A0(n7306));
   OAI21X1TS U870 (.Y(n3935), 
	.B0(n7316), 
	.A1(n3933), 
	.A0(n7311));
   OAI21X1TS U1014 (.Y(n4110), 
	.B0(n7425), 
	.A1(n4108), 
	.A0(n7420));
   AOI21X1TS U1013 (.Y(n5553), 
	.B0(FE_OFN811_n7619), 
	.A1(n4110), 
	.A0(\fifo_to_fir/fifo_cell5/controller/valid_read ));
   OAI21X1TS U1024 (.Y(n4120), 
	.B0(n4122), 
	.A1(n4118), 
	.A0(n7435));
   OAI21X1TS U1021 (.Y(n5558), 
	.B0(n4120), 
	.A1(n4119), 
	.A0(\fifo_to_fir/fifo_cell3/data_out/N35 ));
   OAI211X1TS U1067 (.Y(n4174), 
	.C0(n9473), 
	.B0(\fifo_to_fir/hang[1] ), 
	.A1(n4176), 
	.A0(n8791));
   AOI21X1TS U884 (.Y(n5510), 
	.B0(FE_OFN794_n7619), 
	.A1(n3950), 
	.A0(\fifo_to_fft/fifo_cell2/controller/valid_read ));
   AOI21X1TS U1028 (.Y(n5562), 
	.B0(FE_OFN784_n7619), 
	.A1(n4125), 
	.A0(\fifo_to_fir/fifo_cell2/controller/valid_read ));
   OAI21X1TS U882 (.Y(n5509), 
	.B0(n3950), 
	.A1(n3949), 
	.A0(\fifo_to_fft/fifo_cell2/data_out/N35 ));
   OAI21X1TS U1026 (.Y(n5561), 
	.B0(n4125), 
	.A1(n4124), 
	.A0(\fifo_to_fir/fifo_cell2/data_out/N35 ));
   NOR2X1TS U800 (.Y(n3826), 
	.B(n7610), 
	.A(FE_OFN973_n7207));
   OAI21X1TS U787 (.Y(n5459), 
	.B0(n3824), 
	.A1(n3823), 
	.A0(n7610));
   NOR2X1TS U2737 (.Y(n4841), 
	.B(n4840), 
	.A(instruction[2]));
   NOR2X1TS U2733 (.Y(n3848), 
	.B(n4840), 
	.A(n3455));
   AOI32X1TS U2731 (.Y(n4449), 
	.B1(n9463), 
	.B0(n4456), 
	.A2(n3710), 
	.A1(n9464), 
	.A0(\router/iir_write_done ));
   NOR2X1TS U1434 (.Y(n4452), 
	.B(n4456), 
	.A(n3710));
   AOI32X1TS U1430 (.Y(n4451), 
	.B1(n9464), 
	.B0(n4453), 
	.A2(n4452), 
	.A1(n9464), 
	.A0(\router/iir_write_done ));
   OAI31X1TS U1429 (.Y(n5703), 
	.B0(n4451), 
	.A2(n4450), 
	.A1(n4449), 
	.A0(n4204));
   NOR2X1TS U3442 (.Y(\fifo_to_fir/fifo_cell0/N7 ), 
	.B(n7445), 
	.A(\fifo_to_fir/fifo_cell0/control_signal ));
   NOR2X1TS U3586 (.Y(\fifo_to_fft/fifo_cell0/N7 ), 
	.B(n7336), 
	.A(\fifo_to_fft/fifo_cell0/control_signal ));
   NAND2X1TS U3855 (.Y(n4506), 
	.B(\fifo_from_fft/fifo_cell12/reg_gtok/token ), 
	.A(FE_OFN722_n4643));
   NAND2X1TS U3869 (.Y(n4578), 
	.B(\fifo_from_fft/fifo_cell0/reg_gtok/token ), 
	.A(FE_OFN720_n4643));
   INVX2TS U3380 (.Y(n4176), 
	.A(n4030));
   NOR3X1TS U3378 (.Y(n5203), 
	.C(\fifo_to_fir/fifo_cell3/controller/valid_read ), 
	.B(\fifo_to_fir/fifo_cell3/controller/write_enable ), 
	.A(n7435));
   NOR3X1TS U3374 (.Y(n5202), 
	.C(\fifo_to_fir/fifo_cell4/controller/valid_read ), 
	.B(\fifo_to_fir/fifo_cell4/controller/write_enable ), 
	.A(n7430));
   INVX2TS U3372 (.Y(n4170), 
	.A(n4034));
   INVX2TS U3364 (.Y(n4164), 
	.A(n4038));
   INVX2TS U3360 (.Y(n4161), 
	.A(n4040));
   INVX2TS U3352 (.Y(n4155), 
	.A(n4044));
   INVX2TS U3348 (.Y(n4152), 
	.A(n4046));
   NOR3X1TS U3338 (.Y(n5193), 
	.C(\fifo_to_fir/fifo_cell13/controller/valid_read ), 
	.B(\fifo_to_fir/fifo_cell13/controller/write_enable ), 
	.A(n7361));
   INVX2TS U3336 (.Y(n4143), 
	.A(n4052));
   INVX2TS U3332 (.Y(n4140), 
	.A(n4054));
   NOR3X1TS U3525 (.Y(n5246), 
	.C(\fifo_to_fft/fifo_cell2/controller/valid_read ), 
	.B(\fifo_to_fft/fifo_cell2/controller/write_enable ), 
	.A(n7331));
   AOI31X1TS U3524 (.Y(n3855), 
	.B0(\fifo_to_fft/hold[2] ), 
	.A2(n5246), 
	.A1(\fifo_to_fft/fifo_cell2/data_out/N35 ), 
	.A0(n3952));
   INVX2TS U3515 (.Y(n3995), 
	.A(n3859));
   INVX2TS U3507 (.Y(n3989), 
	.A(n3863));
   INVX2TS U3503 (.Y(n3986), 
	.A(n3865));
   INVX2TS U3495 (.Y(n3980), 
	.A(n3869));
   INVX2TS U3491 (.Y(n3977), 
	.A(n3871));
   INVX2TS U3475 (.Y(n3965), 
	.A(n3879));
   NOR2X1TS U1920 (.Y(n4562), 
	.B(FE_OFN314_n4561), 
	.A(FE_OFN835_n7619));
   NOR2X1TS U2551 (.Y(n4748), 
	.B(FE_OFN658_n4747), 
	.A(FE_OFN846_n7619));
   NOR2X1TS U2588 (.Y(n4754), 
	.B(n8137), 
	.A(FE_OFN833_n7619));
   NOR2X1TS U1957 (.Y(n4568), 
	.B(n8472), 
	.A(FE_OFN835_n7619));
   NOR2X1TS U1994 (.Y(n4574), 
	.B(FE_OFN337_n4573), 
	.A(FE_OFN840_n7619));
   NOR2X1TS U2625 (.Y(n4760), 
	.B(FE_OFN672_n4759), 
	.A(FE_OFN841_n7619));
   NOR4XLTS U2722 (.Y(n3834), 
	.D(\router/iir_get_req_reg ), 
	.C(FE_OFN1284_router_ram_read_enable_reg), 
	.B(\router/fir_get_req_reg ), 
	.A(FE_OFN1282_router_fft_get_req_reg));
   INVX2TS U2703 (.Y(n3828), 
	.A(n3754));
   AOI22XLTS U276 (.Y(n3509), 
	.B1(\router/addr_calc/iir_write_calc/counter/N55 ), 
	.B0(FE_OFN936_n3487), 
	.A1(FE_OFN947_n3486), 
	.A0(\router/addr_calc/iir_write_calc/count[9] ));
   OAI32XLTS U608 (.Y(n3706), 
	.B1(FE_OFN977_n9462), 
	.B0(\router/fft_read_done ), 
	.A2(n3709), 
	.A1(n3708), 
	.A0(n9432));
   OAI21X1TS U885 (.Y(n3950), 
	.B0(n3952), 
	.A1(n3948), 
	.A0(n7331));
   OAI21X1TS U1029 (.Y(n4125), 
	.B0(n4127), 
	.A1(n4123), 
	.A0(n7440));
   NOR2XLTS U2729 (.Y(n4830), 
	.B(\router/ram_read_enable_reg ), 
	.A(\router/fft_get_req_reg ));
   AOI21XLTS U1439 (.Y(n4204), 
	.B0(n4200), 
	.A1(n7211), 
	.A0(\router/fir_write_done ));
   OAI31X1TS U1103 (.Y(n5573), 
	.B0(n4201), 
	.A2(n4200), 
	.A1(\router/fir_write_done ), 
	.A0(FE_OFN843_n7619));
   OAI211X1TS U225 (.Y(\router/data_cntl/N134 ), 
	.C0(n3481), 
	.B0(n3480), 
	.A1(n3479), 
	.A0(\router/data_cntl/fft_full_flag ));
   NAND2X1TS U3712 (.Y(n4692), 
	.B(\fifo_from_fir/fifo_cell12/reg_gtok/token ), 
	.A(FE_OFN735_n4829));
   NOR2X1TS U1550 (.Y(n4502), 
	.B(n8711), 
	.A(FE_OFN847_n7619));
   NOR2X1TS U2181 (.Y(n4688), 
	.B(n8376), 
	.A(FE_OFN828_n7619));
   NOR2X1TS U1661 (.Y(n4520), 
	.B(FE_OFN210_n4519), 
	.A(FE_OFN836_n7619));
   NAND2X1TS U2715 (.Y(n4644), 
	.B(n7606), 
	.A(FE_OFN776_n3829));
   NAND2X1TS U2073 (.Y(n3755), 
	.B(FE_OFN776_n3829), 
	.A(n9435));
   AOI22XLTS U274 (.Y(n3508), 
	.B1(\router/addr_calc/iir_write_calc/counter/N56 ), 
	.B0(FE_OFN936_n3487), 
	.A1(FE_OFN948_n3486), 
	.A0(n7104));
   AOI22XLTS U270 (.Y(n3506), 
	.B1(\router/addr_calc/iir_write_calc/counter/N58 ), 
	.B0(FE_OFN935_n3487), 
	.A1(FE_OFN948_n3486), 
	.A0(n7115));
   AOI211X1TS U789 (.Y(n3823), 
	.C0(n3828), 
	.B0(n3827), 
	.A1(n7608), 
	.A0(n3826));
   NOR3X1TS U3757 (.Y(n5312), 
	.C(\fifo_from_fft/fifo_cell15/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell15/controller/write_enable ), 
	.A(n7455));
   AOI32X1TS U2714 (.Y(n3832), 
	.B1(FE_OFN776_n3829), 
	.B0(n9433), 
	.A2(n9389), 
	.A1(FE_OFN776_n3829), 
	.A0(FE_OFN990_n9431));
   AOI211X1TS U229 (.Y(\router/data_cntl/N135 ), 
	.C0(n3483), 
	.B0(FE_OFN979_n9462), 
	.A1(FE_OFN1217_n3478), 
	.A0(n3482));
   AOI211X1TS U220 (.Y(\router/data_cntl/N137 ), 
	.C0(n3473), 
	.B0(FE_OFN973_n7207), 
	.A1(n3467), 
	.A0(n3471));
   AOI211X1TS U611 (.Y(n3705), 
	.C0(n3715), 
	.B0(n3714), 
	.A1(n3713), 
	.A0(n3712));
   NOR2X4TS U610 (.Y(ram_read_enable), 
	.B(n7610), 
	.A(n3705));
   ADDHXLTS \add_x_22_5/U1_1_27  (.S(\router/addr_calc/iir_write_calc/counter/N73 ), 
	.CO(\add_x_22_5/carry[28] ), 
	.B(\add_x_22_5/carry[27] ), 
	.A(FE_OFN1439_router_addr_calc_iir_write_calc_count_27_));
   ADDHXLTS \add_x_22_5/U1_1_26  (.S(\router/addr_calc/iir_write_calc/counter/N72 ), 
	.CO(\add_x_22_5/carry[27] ), 
	.B(\add_x_22_5/carry[26] ), 
	.A(n7181));
   ADDHXLTS \add_x_22_5/U1_1_25  (.S(\router/addr_calc/iir_write_calc/counter/N71 ), 
	.CO(\add_x_22_5/carry[26] ), 
	.B(\add_x_22_5/carry[25] ), 
	.A(n7175));
   ADDHXLTS \add_x_22_5/U1_1_24  (.S(\router/addr_calc/iir_write_calc/counter/N70 ), 
	.CO(\add_x_22_5/carry[25] ), 
	.B(\add_x_22_5/carry[24] ), 
	.A(n7169));
   ADDHXLTS \add_x_22_5/U1_1_23  (.S(\router/addr_calc/iir_write_calc/counter/N69 ), 
	.CO(\add_x_22_5/carry[24] ), 
	.B(\add_x_22_5/carry[23] ), 
	.A(FE_OFN1244_router_addr_calc_iir_write_calc_count_23_));
   ADDHXLTS \add_x_22_5/U1_1_22  (.S(\router/addr_calc/iir_write_calc/counter/N68 ), 
	.CO(\add_x_22_5/carry[23] ), 
	.B(\add_x_22_5/carry[22] ), 
	.A(n7163));
   ADDHXLTS \add_x_22_5/U1_1_21  (.S(\router/addr_calc/iir_write_calc/counter/N67 ), 
	.CO(\add_x_22_5/carry[22] ), 
	.B(\add_x_22_5/carry[21] ), 
	.A(n7156));
   ADDHXLTS \add_x_22_5/U1_1_20  (.S(\router/addr_calc/iir_write_calc/counter/N66 ), 
	.CO(\add_x_22_5/carry[21] ), 
	.B(\add_x_22_5/carry[20] ), 
	.A(n7150));
   ADDHXLTS \add_x_22_5/U1_1_19  (.S(\router/addr_calc/iir_write_calc/counter/N65 ), 
	.CO(\add_x_22_5/carry[20] ), 
	.B(\add_x_22_5/carry[19] ), 
	.A(FE_OFN1440_router_addr_calc_iir_write_calc_count_19_));
   ADDHXLTS \add_x_22_5/U1_1_18  (.S(\router/addr_calc/iir_write_calc/counter/N64 ), 
	.CO(\add_x_22_5/carry[19] ), 
	.B(\add_x_22_5/carry[18] ), 
	.A(n7144));
   ADDHXLTS \add_x_22_5/U1_1_17  (.S(\router/addr_calc/iir_write_calc/counter/N63 ), 
	.CO(\add_x_22_5/carry[18] ), 
	.B(\add_x_22_5/carry[17] ), 
	.A(n7138));
   ADDHXLTS \add_x_22_5/U1_1_16  (.S(\router/addr_calc/iir_write_calc/counter/N62 ), 
	.CO(\add_x_22_5/carry[17] ), 
	.B(\add_x_22_5/carry[16] ), 
	.A(FE_OFN1441_router_addr_calc_iir_write_calc_count_16_));
   ADDHXLTS \add_x_22_5/U1_1_15  (.S(\router/addr_calc/iir_write_calc/counter/N61 ), 
	.CO(\add_x_22_5/carry[16] ), 
	.B(\add_x_22_5/carry[15] ), 
	.A(n7132));
   ADDHXLTS \add_x_22_5/U1_1_14  (.S(\router/addr_calc/iir_write_calc/counter/N60 ), 
	.CO(\add_x_22_5/carry[15] ), 
	.B(\add_x_22_5/carry[14] ), 
	.A(n7126));
   ADDHXLTS \add_x_22_5/U1_1_13  (.S(\router/addr_calc/iir_write_calc/counter/N59 ), 
	.CO(\add_x_22_5/carry[14] ), 
	.B(\add_x_22_5/carry[13] ), 
	.A(n7121));
   ADDHXLTS \add_x_22_5/U1_1_12  (.S(\router/addr_calc/iir_write_calc/counter/N58 ), 
	.CO(\add_x_22_5/carry[13] ), 
	.B(\add_x_22_5/carry[12] ), 
	.A(n7115));
   ADDHXLTS \add_x_22_5/U1_1_11  (.S(\router/addr_calc/iir_write_calc/counter/N57 ), 
	.CO(\add_x_22_5/carry[12] ), 
	.B(\add_x_22_5/carry[11] ), 
	.A(n7109));
   ADDHXLTS \add_x_22_5/U1_1_10  (.S(\router/addr_calc/iir_write_calc/counter/N56 ), 
	.CO(\add_x_22_5/carry[11] ), 
	.B(\add_x_22_5/carry[10] ), 
	.A(n7104));
   ADDHXLTS \add_x_22_5/U1_1_9  (.S(\router/addr_calc/iir_write_calc/counter/N55 ), 
	.CO(\add_x_22_5/carry[10] ), 
	.B(\add_x_22_5/carry[9] ), 
	.A(FE_OFN1280_router_addr_calc_iir_write_calc_count_9_));
   ADDHXLTS \add_x_22_5/U1_1_8  (.S(\router/addr_calc/iir_write_calc/counter/N54 ), 
	.CO(\add_x_22_5/carry[9] ), 
	.B(\add_x_22_5/carry[8] ), 
	.A(n7098));
   ADDHXLTS \add_x_22_5/U1_1_7  (.S(\router/addr_calc/iir_write_calc/counter/N53 ), 
	.CO(\add_x_22_5/carry[8] ), 
	.B(\add_x_22_5/carry[7] ), 
	.A(n7092));
   ADDHXLTS \add_x_22_5/U1_1_6  (.S(\router/addr_calc/iir_write_calc/counter/N52 ), 
	.CO(\add_x_22_5/carry[7] ), 
	.B(\add_x_22_5/carry[6] ), 
	.A(n7089));
   ADDHXLTS \add_x_22_5/U1_1_5  (.S(\router/addr_calc/iir_write_calc/counter/N51 ), 
	.CO(\add_x_22_5/carry[6] ), 
	.B(\add_x_22_5/carry[5] ), 
	.A(FE_OFN1281_router_addr_calc_iir_write_calc_count_5_));
   ADDHXLTS \add_x_22_5/U1_1_4  (.S(\router/addr_calc/iir_write_calc/counter/N50 ), 
	.CO(\add_x_22_5/carry[5] ), 
	.B(\add_x_22_5/carry[4] ), 
	.A(n7095));
   ADDHXLTS \add_x_22_5/U1_1_3  (.S(\router/addr_calc/iir_write_calc/counter/N49 ), 
	.CO(\add_x_22_5/carry[4] ), 
	.B(\add_x_22_5/carry[3] ), 
	.A(n7101));
   ADDHXLTS \add_x_22_5/U1_1_2  (.S(\router/addr_calc/iir_write_calc/counter/N48 ), 
	.CO(\add_x_22_5/carry[3] ), 
	.B(\add_x_22_5/carry[2] ), 
	.A(FE_OFN1825_n7107));
   ADDHXLTS \add_x_22_5/U1_1_1  (.S(\router/addr_calc/iir_write_calc/counter/N47 ), 
	.CO(\add_x_22_5/carry[2] ), 
	.B(FE_OFN1442_router_addr_calc_iir_write_calc_count_0_), 
	.A(n7112));
   ADDHXLTS \add_x_22_3/U1_1_27  (.S(\router/addr_calc/fir_write_calc/counter/N73 ), 
	.CO(\add_x_22_3/carry[28] ), 
	.B(\add_x_22_3/carry[27] ), 
	.A(\router/addr_calc/fir_write_calc/count[27] ));
   ADDHXLTS \add_x_22_3/U1_1_26  (.S(\router/addr_calc/fir_write_calc/counter/N72 ), 
	.CO(\add_x_22_3/carry[27] ), 
	.B(\add_x_22_3/carry[26] ), 
	.A(n7136));
   ADDHXLTS \add_x_22_3/U1_1_25  (.S(\router/addr_calc/fir_write_calc/counter/N71 ), 
	.CO(\add_x_22_3/carry[26] ), 
	.B(\add_x_22_3/carry[25] ), 
	.A(n7142));
   ADDHXLTS \add_x_22_3/U1_1_24  (.S(\router/addr_calc/fir_write_calc/counter/N70 ), 
	.CO(\add_x_22_3/carry[25] ), 
	.B(\add_x_22_3/carry[24] ), 
	.A(n7148));
   ADDHXLTS \add_x_22_3/U1_1_23  (.S(\router/addr_calc/fir_write_calc/counter/N69 ), 
	.CO(\add_x_22_3/carry[24] ), 
	.B(\add_x_22_3/carry[23] ), 
	.A(FE_OFN1248_router_addr_calc_fir_write_calc_count_23_));
   ADDHXLTS \add_x_22_3/U1_1_22  (.S(\router/addr_calc/fir_write_calc/counter/N68 ), 
	.CO(\add_x_22_3/carry[23] ), 
	.B(\add_x_22_3/carry[22] ), 
	.A(n7154));
   ADDHXLTS \add_x_22_3/U1_1_21  (.S(\router/addr_calc/fir_write_calc/counter/N67 ), 
	.CO(\add_x_22_3/carry[22] ), 
	.B(\add_x_22_3/carry[21] ), 
	.A(n7160));
   ADDHXLTS \add_x_22_3/U1_1_20  (.S(\router/addr_calc/fir_write_calc/counter/N66 ), 
	.CO(\add_x_22_3/carry[21] ), 
	.B(\add_x_22_3/carry[20] ), 
	.A(FE_OFN1257_n7165));
   ADDHXLTS \add_x_22_3/U1_1_19  (.S(\router/addr_calc/fir_write_calc/counter/N65 ), 
	.CO(\add_x_22_3/carry[20] ), 
	.B(\add_x_22_3/carry[19] ), 
	.A(\router/addr_calc/fir_write_calc/count[19] ));
   ADDHXLTS \add_x_22_3/U1_1_18  (.S(\router/addr_calc/fir_write_calc/counter/N64 ), 
	.CO(\add_x_22_3/carry[19] ), 
	.B(\add_x_22_3/carry[18] ), 
	.A(n7171));
   ADDHXLTS \add_x_22_3/U1_1_17  (.S(\router/addr_calc/fir_write_calc/counter/N63 ), 
	.CO(\add_x_22_3/carry[18] ), 
	.B(\add_x_22_3/carry[17] ), 
	.A(n7177));
   ADDHXLTS \add_x_22_3/U1_1_16  (.S(\router/addr_calc/fir_write_calc/counter/N62 ), 
	.CO(\add_x_22_3/carry[17] ), 
	.B(\add_x_22_3/carry[16] ), 
	.A(\router/addr_calc/fir_write_calc/count[16] ));
   ADDHXLTS \add_x_22_3/U1_1_15  (.S(\router/addr_calc/fir_write_calc/counter/N61 ), 
	.CO(\add_x_22_3/carry[16] ), 
	.B(\add_x_22_3/carry[15] ), 
	.A(n7183));
   ADDHXLTS \add_x_22_3/U1_1_14  (.S(\router/addr_calc/fir_write_calc/counter/N60 ), 
	.CO(\add_x_22_3/carry[15] ), 
	.B(\add_x_22_3/carry[14] ), 
	.A(n7189));
   ADDHXLTS \add_x_22_3/U1_1_13  (.S(\router/addr_calc/fir_write_calc/counter/N59 ), 
	.CO(\add_x_22_3/carry[14] ), 
	.B(\add_x_22_3/carry[13] ), 
	.A(n7195));
   ADDHXLTS \add_x_22_3/U1_1_12  (.S(\router/addr_calc/fir_write_calc/counter/N58 ), 
	.CO(\add_x_22_3/carry[13] ), 
	.B(\add_x_22_3/carry[12] ), 
	.A(n7201));
   ADDHXLTS \add_x_22_3/U1_1_11  (.S(\router/addr_calc/fir_write_calc/counter/N57 ), 
	.CO(\add_x_22_3/carry[12] ), 
	.B(\add_x_22_3/carry[11] ), 
	.A(n7205));
   ADDHXLTS \add_x_22_3/U1_1_10  (.S(\router/addr_calc/fir_write_calc/counter/N56 ), 
	.CO(\add_x_22_3/carry[11] ), 
	.B(\add_x_22_3/carry[10] ), 
	.A(n7209));
   ADDHXLTS \add_x_22_3/U1_1_9  (.S(\router/addr_calc/fir_write_calc/counter/N55 ), 
	.CO(\add_x_22_3/carry[10] ), 
	.B(\add_x_22_3/carry[9] ), 
	.A(FE_OFN1266_router_addr_calc_fir_write_calc_count_9_));
   ADDHXLTS \add_x_22_3/U1_1_8  (.S(\router/addr_calc/fir_write_calc/counter/N54 ), 
	.CO(\add_x_22_3/carry[9] ), 
	.B(\add_x_22_3/carry[8] ), 
	.A(n7214));
   ADDHXLTS \add_x_22_3/U1_1_7  (.S(\router/addr_calc/fir_write_calc/counter/N53 ), 
	.CO(\add_x_22_3/carry[8] ), 
	.B(\add_x_22_3/carry[7] ), 
	.A(n7219));
   ADDHXLTS \add_x_22_3/U1_1_6  (.S(\router/addr_calc/fir_write_calc/counter/N52 ), 
	.CO(\add_x_22_3/carry[7] ), 
	.B(\add_x_22_3/carry[6] ), 
	.A(n7224));
   ADDHXLTS \add_x_22_3/U1_1_5  (.S(\router/addr_calc/fir_write_calc/counter/N51 ), 
	.CO(\add_x_22_3/carry[6] ), 
	.B(\add_x_22_3/carry[5] ), 
	.A(FE_OFN1272_router_addr_calc_fir_write_calc_count_5_));
   ADDHXLTS \add_x_22_3/U1_1_4  (.S(\router/addr_calc/fir_write_calc/counter/N50 ), 
	.CO(\add_x_22_3/carry[5] ), 
	.B(\add_x_22_3/carry[4] ), 
	.A(n7229));
   ADDHXLTS \add_x_22_3/U1_1_3  (.S(\router/addr_calc/fir_write_calc/counter/N49 ), 
	.CO(\add_x_22_3/carry[4] ), 
	.B(\add_x_22_3/carry[3] ), 
	.A(n7234));
   ADDHXLTS \add_x_22_3/U1_1_2  (.S(\router/addr_calc/fir_write_calc/counter/N48 ), 
	.CO(\add_x_22_3/carry[3] ), 
	.B(\add_x_22_3/carry[2] ), 
	.A(n7239));
   ADDHXLTS \add_x_22_2/U1_1_27  (.S(\router/addr_calc/fir_read_calc/counter/N73 ), 
	.CO(\add_x_22_2/carry[28] ), 
	.B(\add_x_22_2/carry[27] ), 
	.A(FE_OFN1239_router_addr_calc_fir_read_calc_count_27_));
   ADDHXLTS \add_x_22_2/U1_1_26  (.S(\router/addr_calc/fir_read_calc/counter/N72 ), 
	.CO(\add_x_22_2/carry[27] ), 
	.B(\add_x_22_2/carry[26] ), 
	.A(FE_OFN1241_n7264));
   ADDHXLTS \add_x_22_2/U1_1_25  (.S(\router/addr_calc/fir_read_calc/counter/N71 ), 
	.CO(\add_x_22_2/carry[26] ), 
	.B(\add_x_22_2/carry[25] ), 
	.A(n7269));
   ADDHXLTS \add_x_22_2/U1_1_24  (.S(\router/addr_calc/fir_read_calc/counter/N70 ), 
	.CO(\add_x_22_2/carry[25] ), 
	.B(\add_x_22_2/carry[24] ), 
	.A(n7274));
   ADDHXLTS \add_x_22_2/U1_1_23  (.S(\router/addr_calc/fir_read_calc/counter/N69 ), 
	.CO(\add_x_22_2/carry[24] ), 
	.B(\add_x_22_2/carry[23] ), 
	.A(FE_OFN1247_router_addr_calc_fir_read_calc_count_23_));
   ADDHXLTS \add_x_22_2/U1_1_22  (.S(\router/addr_calc/fir_read_calc/counter/N68 ), 
	.CO(\add_x_22_2/carry[23] ), 
	.B(\add_x_22_2/carry[22] ), 
	.A(n7279));
   ADDHXLTS \add_x_22_2/U1_1_21  (.S(\router/addr_calc/fir_read_calc/counter/N67 ), 
	.CO(\add_x_22_2/carry[22] ), 
	.B(\add_x_22_2/carry[21] ), 
	.A(n7284));
   ADDHXLTS \add_x_22_2/U1_1_20  (.S(\router/addr_calc/fir_read_calc/counter/N66 ), 
	.CO(\add_x_22_2/carry[21] ), 
	.B(\add_x_22_2/carry[20] ), 
	.A(FE_OFN1256_n7288));
   ADDHXLTS \add_x_22_2/U1_1_19  (.S(\router/addr_calc/fir_read_calc/counter/N65 ), 
	.CO(\add_x_22_2/carry[20] ), 
	.B(\add_x_22_2/carry[19] ), 
	.A(\router/addr_calc/fir_read_calc/count[19] ));
   ADDHXLTS \add_x_22_2/U1_1_18  (.S(\router/addr_calc/fir_read_calc/counter/N64 ), 
	.CO(\add_x_22_2/carry[19] ), 
	.B(\add_x_22_2/carry[18] ), 
	.A(n7293));
   ADDHXLTS \add_x_22_2/U1_1_17  (.S(\router/addr_calc/fir_read_calc/counter/N63 ), 
	.CO(\add_x_22_2/carry[18] ), 
	.B(\add_x_22_2/carry[17] ), 
	.A(FE_OFN1262_n7298));
   ADDHXLTS \add_x_22_2/U1_1_16  (.S(\router/addr_calc/fir_read_calc/counter/N62 ), 
	.CO(\add_x_22_2/carry[17] ), 
	.B(\add_x_22_2/carry[16] ), 
	.A(FE_OFN1265_n7303));
   ADDHXLTS \add_x_22_2/U1_1_15  (.S(\router/addr_calc/fir_read_calc/counter/N61 ), 
	.CO(\add_x_22_2/carry[16] ), 
	.B(\add_x_22_2/carry[15] ), 
	.A(FE_OFN1271_router_addr_calc_fir_read_calc_count_15_));
   ADDHXLTS \add_x_22_2/U1_1_14  (.S(\router/addr_calc/fir_read_calc/counter/N60 ), 
	.CO(\add_x_22_2/carry[15] ), 
	.B(\add_x_22_2/carry[14] ), 
	.A(FE_OFN1277_n7308));
   ADDHXLTS \add_x_22_2/U1_1_13  (.S(\router/addr_calc/fir_read_calc/counter/N59 ), 
	.CO(\add_x_22_2/carry[14] ), 
	.B(\add_x_22_2/carry[13] ), 
	.A(n7313));
   ADDHXLTS \add_x_22_2/U1_1_12  (.S(\router/addr_calc/fir_read_calc/counter/N58 ), 
	.CO(\add_x_22_2/carry[13] ), 
	.B(\add_x_22_2/carry[12] ), 
	.A(n7318));
   ADDHXLTS \add_x_22_2/U1_1_11  (.S(\router/addr_calc/fir_read_calc/counter/N57 ), 
	.CO(\add_x_22_2/carry[12] ), 
	.B(\add_x_22_2/carry[11] ), 
	.A(n7323));
   ADDHXLTS \add_x_22_2/U1_1_10  (.S(\router/addr_calc/fir_read_calc/counter/N56 ), 
	.CO(\add_x_22_2/carry[11] ), 
	.B(\add_x_22_2/carry[10] ), 
	.A(FE_OFN1279_n7328));
   ADDHXLTS \add_x_22_2/U1_1_9  (.S(\router/addr_calc/fir_read_calc/counter/N55 ), 
	.CO(\add_x_22_2/carry[10] ), 
	.B(\add_x_22_2/carry[9] ), 
	.A(FE_OFN1269_router_addr_calc_fir_read_calc_count_9_));
   ADDHXLTS \add_x_22_2/U1_1_8  (.S(\router/addr_calc/fir_read_calc/counter/N54 ), 
	.CO(\add_x_22_2/carry[9] ), 
	.B(\add_x_22_2/carry[8] ), 
	.A(FE_OFN1278_n7333));
   ADDHXLTS \add_x_22_2/U1_1_7  (.S(\router/addr_calc/fir_read_calc/counter/N53 ), 
	.CO(\add_x_22_2/carry[8] ), 
	.B(\add_x_22_2/carry[7] ), 
	.A(n7338));
   ADDHXLTS \add_x_22_2/U1_1_6  (.S(\router/addr_calc/fir_read_calc/counter/N52 ), 
	.CO(\add_x_22_2/carry[7] ), 
	.B(\add_x_22_2/carry[6] ), 
	.A(n7343));
   ADDHXLTS \add_x_22_2/U1_1_5  (.S(\router/addr_calc/fir_read_calc/counter/N51 ), 
	.CO(\add_x_22_2/carry[6] ), 
	.B(\add_x_22_2/carry[5] ), 
	.A(FE_OFN1824_router_addr_calc_fir_read_calc_count_5_));
   ADDHXLTS \add_x_22_2/U1_1_4  (.S(\router/addr_calc/fir_read_calc/counter/N50 ), 
	.CO(\add_x_22_2/carry[5] ), 
	.B(\add_x_22_2/carry[4] ), 
	.A(n7348));
   ADDHXLTS \add_x_22_2/U1_1_3  (.S(\router/addr_calc/fir_read_calc/counter/N49 ), 
	.CO(\add_x_22_2/carry[4] ), 
	.B(\add_x_22_2/carry[3] ), 
	.A(FE_OFN1275_n7353));
   ADDHXLTS \add_x_22_2/U1_1_2  (.S(\router/addr_calc/fir_read_calc/counter/N48 ), 
	.CO(\add_x_22_2/carry[3] ), 
	.B(\add_x_22_2/carry[2] ), 
	.A(FE_OFN1274_n7358));
   ADDHXLTS \add_x_22_1/U1_1_29  (.S(\router/addr_calc/fft_write_calc/counter/N75 ), 
	.CO(\add_x_22_1/carry[30] ), 
	.B(\add_x_22_1/carry[29] ), 
	.A(FE_OFN1233_router_addr_calc_fft_write_calc_count_29_));
   ADDHXLTS \add_x_22_1/U1_1_27  (.S(\router/addr_calc/fft_write_calc/counter/N73 ), 
	.CO(\add_x_22_1/carry[28] ), 
	.B(\add_x_22_1/carry[27] ), 
	.A(FE_OFN1238_router_addr_calc_fft_write_calc_count_27_));
   ADDHXLTS \add_x_22_1/U1_1_26  (.S(\router/addr_calc/fft_write_calc/counter/N72 ), 
	.CO(\add_x_22_1/carry[27] ), 
	.B(\add_x_22_1/carry[26] ), 
	.A(n7378));
   ADDHXLTS \add_x_22_1/U1_1_25  (.S(\router/addr_calc/fft_write_calc/counter/N71 ), 
	.CO(\add_x_22_1/carry[26] ), 
	.B(\add_x_22_1/carry[25] ), 
	.A(n7383));
   ADDHXLTS \add_x_22_1/U1_1_24  (.S(\router/addr_calc/fft_write_calc/counter/N70 ), 
	.CO(\add_x_22_1/carry[25] ), 
	.B(\add_x_22_1/carry[24] ), 
	.A(n7388));
   ADDHXLTS \add_x_22_1/U1_1_23  (.S(\router/addr_calc/fft_write_calc/counter/N69 ), 
	.CO(\add_x_22_1/carry[24] ), 
	.B(\add_x_22_1/carry[23] ), 
	.A(FE_OFN1246_router_addr_calc_fft_write_calc_count_23_));
   ADDHXLTS \add_x_22_1/U1_1_22  (.S(\router/addr_calc/fft_write_calc/counter/N68 ), 
	.CO(\add_x_22_1/carry[23] ), 
	.B(\add_x_22_1/carry[22] ), 
	.A(n7393));
   ADDHXLTS \add_x_22_1/U1_1_21  (.S(\router/addr_calc/fft_write_calc/counter/N67 ), 
	.CO(\add_x_22_1/carry[22] ), 
	.B(\add_x_22_1/carry[21] ), 
	.A(n7398));
   ADDHXLTS \add_x_22_1/U1_1_20  (.S(\router/addr_calc/fft_write_calc/counter/N66 ), 
	.CO(\add_x_22_1/carry[21] ), 
	.B(\add_x_22_1/carry[20] ), 
	.A(FE_OFN1255_n7402));
   ADDHXLTS \add_x_22_1/U1_1_19  (.S(\router/addr_calc/fft_write_calc/counter/N65 ), 
	.CO(\add_x_22_1/carry[20] ), 
	.B(\add_x_22_1/carry[19] ), 
	.A(FE_OFN1259_router_addr_calc_fft_write_calc_count_19_));
   ADDHXLTS \add_x_22_1/U1_1_18  (.S(\router/addr_calc/fft_write_calc/counter/N64 ), 
	.CO(\add_x_22_1/carry[19] ), 
	.B(\add_x_22_1/carry[18] ), 
	.A(n7407));
   ADDHXLTS \add_x_22_1/U1_1_17  (.S(\router/addr_calc/fft_write_calc/counter/N63 ), 
	.CO(\add_x_22_1/carry[18] ), 
	.B(\add_x_22_1/carry[17] ), 
	.A(n7412));
   ADDHXLTS \add_x_22_1/U1_1_16  (.S(\router/addr_calc/fft_write_calc/counter/N62 ), 
	.CO(\add_x_22_1/carry[17] ), 
	.B(\add_x_22_1/carry[16] ), 
	.A(n7417));
   ADDHXLTS \add_x_22_1/U1_1_15  (.S(\router/addr_calc/fft_write_calc/counter/N61 ), 
	.CO(\add_x_22_1/carry[16] ), 
	.B(\add_x_22_1/carry[15] ), 
	.A(FE_OFN1270_router_addr_calc_fft_write_calc_count_15_));
   ADDHXLTS \add_x_22_1/U1_1_14  (.S(\router/addr_calc/fft_write_calc/counter/N60 ), 
	.CO(\add_x_22_1/carry[15] ), 
	.B(\add_x_22_1/carry[14] ), 
	.A(n7422));
   ADDHXLTS \add_x_22_1/U1_1_13  (.S(\router/addr_calc/fft_write_calc/counter/N59 ), 
	.CO(\add_x_22_1/carry[14] ), 
	.B(\add_x_22_1/carry[13] ), 
	.A(n7427));
   ADDHXLTS \add_x_22_1/U1_1_12  (.S(\router/addr_calc/fft_write_calc/counter/N58 ), 
	.CO(\add_x_22_1/carry[13] ), 
	.B(\add_x_22_1/carry[12] ), 
	.A(n7432));
   ADDHXLTS \add_x_22_1/U1_1_11  (.S(\router/addr_calc/fft_write_calc/counter/N57 ), 
	.CO(\add_x_22_1/carry[12] ), 
	.B(\add_x_22_1/carry[11] ), 
	.A(n7437));
   ADDHXLTS \add_x_22_1/U1_1_10  (.S(\router/addr_calc/fft_write_calc/counter/N56 ), 
	.CO(\add_x_22_1/carry[11] ), 
	.B(\add_x_22_1/carry[10] ), 
	.A(n7442));
   ADDHXLTS \add_x_22_1/U1_1_9  (.S(\router/addr_calc/fft_write_calc/counter/N55 ), 
	.CO(\add_x_22_1/carry[10] ), 
	.B(\add_x_22_1/carry[9] ), 
	.A(FE_OFN1268_router_addr_calc_fft_write_calc_count_9_));
   ADDHXLTS \add_x_22_1/U1_1_8  (.S(\router/addr_calc/fft_write_calc/counter/N54 ), 
	.CO(\add_x_22_1/carry[9] ), 
	.B(\add_x_22_1/carry[8] ), 
	.A(n7447));
   ADDHXLTS \add_x_22_1/U1_1_7  (.S(\router/addr_calc/fft_write_calc/counter/N53 ), 
	.CO(\add_x_22_1/carry[8] ), 
	.B(\add_x_22_1/carry[7] ), 
	.A(n7452));
   ADDHXLTS \add_x_22_1/U1_1_6  (.S(\router/addr_calc/fft_write_calc/counter/N52 ), 
	.CO(\add_x_22_1/carry[7] ), 
	.B(\add_x_22_1/carry[6] ), 
	.A(n7457));
   ADDHXLTS \add_x_22_1/U1_1_5  (.S(\router/addr_calc/fft_write_calc/counter/N51 ), 
	.CO(\add_x_22_1/carry[6] ), 
	.B(\add_x_22_1/carry[5] ), 
	.A(n7462));
   ADDHXLTS \add_x_22_1/U1_1_4  (.S(\router/addr_calc/fft_write_calc/counter/N50 ), 
	.CO(\add_x_22_1/carry[5] ), 
	.B(\add_x_22_1/carry[4] ), 
	.A(n7467));
   ADDHXLTS \add_x_22_1/U1_1_3  (.S(\router/addr_calc/fft_write_calc/counter/N49 ), 
	.CO(\add_x_22_1/carry[4] ), 
	.B(\add_x_22_1/carry[3] ), 
	.A(n7472));
   ADDHXLTS \add_x_22_1/U1_1_2  (.S(\router/addr_calc/fft_write_calc/counter/N48 ), 
	.CO(\add_x_22_1/carry[3] ), 
	.B(\add_x_22_1/carry[2] ), 
	.A(n7477));
   ADDHXLTS \add_x_22_0/U1_1_27  (.S(\router/addr_calc/fft_read_calc/counter/N73 ), 
	.CO(\add_x_22_0/carry[28] ), 
	.B(\add_x_22_0/carry[27] ), 
	.A(\router/addr_calc/fft_read_calc/count[27] ));
   ADDHXLTS \add_x_22_0/U1_1_26  (.S(\router/addr_calc/fft_read_calc/counter/N72 ), 
	.CO(\add_x_22_0/carry[27] ), 
	.B(\add_x_22_0/carry[26] ), 
	.A(n7502));
   ADDHXLTS \add_x_22_0/U1_1_25  (.S(\router/addr_calc/fft_read_calc/counter/N71 ), 
	.CO(\add_x_22_0/carry[26] ), 
	.B(\add_x_22_0/carry[25] ), 
	.A(n7507));
   ADDHXLTS \add_x_22_0/U1_1_24  (.S(\router/addr_calc/fft_read_calc/counter/N70 ), 
	.CO(\add_x_22_0/carry[25] ), 
	.B(\add_x_22_0/carry[24] ), 
	.A(n7512));
   ADDHXLTS \add_x_22_0/U1_1_23  (.S(\router/addr_calc/fft_read_calc/counter/N69 ), 
	.CO(\add_x_22_0/carry[24] ), 
	.B(\add_x_22_0/carry[23] ), 
	.A(\router/addr_calc/fft_read_calc/count[23] ));
   ADDHXLTS \add_x_22_0/U1_1_22  (.S(\router/addr_calc/fft_read_calc/counter/N68 ), 
	.CO(\add_x_22_0/carry[23] ), 
	.B(\add_x_22_0/carry[22] ), 
	.A(n7517));
   ADDHXLTS \add_x_22_0/U1_1_21  (.S(\router/addr_calc/fft_read_calc/counter/N67 ), 
	.CO(\add_x_22_0/carry[22] ), 
	.B(\add_x_22_0/carry[21] ), 
	.A(n7522));
   ADDHXLTS \add_x_22_0/U1_1_20  (.S(\router/addr_calc/fft_read_calc/counter/N66 ), 
	.CO(\add_x_22_0/carry[21] ), 
	.B(\add_x_22_0/carry[20] ), 
	.A(n7526));
   ADDHXLTS \add_x_22_0/U1_1_19  (.S(\router/addr_calc/fft_read_calc/counter/N65 ), 
	.CO(\add_x_22_0/carry[20] ), 
	.B(\add_x_22_0/carry[19] ), 
	.A(\router/addr_calc/fft_read_calc/count[19] ));
   ADDHXLTS \add_x_22_0/U1_1_18  (.S(\router/addr_calc/fft_read_calc/counter/N64 ), 
	.CO(\add_x_22_0/carry[19] ), 
	.B(\add_x_22_0/carry[18] ), 
	.A(n7531));
   ADDHXLTS \add_x_22_0/U1_1_17  (.S(\router/addr_calc/fft_read_calc/counter/N63 ), 
	.CO(\add_x_22_0/carry[18] ), 
	.B(\add_x_22_0/carry[17] ), 
	.A(n7536));
   ADDHXLTS \add_x_22_0/U1_1_16  (.S(\router/addr_calc/fft_read_calc/counter/N62 ), 
	.CO(\add_x_22_0/carry[17] ), 
	.B(\add_x_22_0/carry[16] ), 
	.A(FE_OFN1263_router_addr_calc_fft_read_calc_count_16_));
   ADDHXLTS \add_x_22_0/U1_1_15  (.S(\router/addr_calc/fft_read_calc/counter/N61 ), 
	.CO(\add_x_22_0/carry[16] ), 
	.B(\add_x_22_0/carry[15] ), 
	.A(n7541));
   ADDHXLTS \add_x_22_0/U1_1_14  (.S(\router/addr_calc/fft_read_calc/counter/N60 ), 
	.CO(\add_x_22_0/carry[15] ), 
	.B(\add_x_22_0/carry[14] ), 
	.A(n7546));
   ADDHXLTS \add_x_22_0/U1_1_13  (.S(\router/addr_calc/fft_read_calc/counter/N59 ), 
	.CO(\add_x_22_0/carry[14] ), 
	.B(\add_x_22_0/carry[13] ), 
	.A(n7551));
   ADDHXLTS \add_x_22_0/U1_1_12  (.S(\router/addr_calc/fft_read_calc/counter/N58 ), 
	.CO(\add_x_22_0/carry[13] ), 
	.B(\add_x_22_0/carry[12] ), 
	.A(n7556));
   ADDHXLTS \add_x_22_0/U1_1_11  (.S(\router/addr_calc/fft_read_calc/counter/N57 ), 
	.CO(\add_x_22_0/carry[12] ), 
	.B(\add_x_22_0/carry[11] ), 
	.A(n7561));
   ADDHXLTS \add_x_22_0/U1_1_10  (.S(\router/addr_calc/fft_read_calc/counter/N56 ), 
	.CO(\add_x_22_0/carry[11] ), 
	.B(\add_x_22_0/carry[10] ), 
	.A(n7566));
   ADDHXLTS \add_x_22_0/U1_1_9  (.S(\router/addr_calc/fft_read_calc/counter/N55 ), 
	.CO(\add_x_22_0/carry[10] ), 
	.B(\add_x_22_0/carry[9] ), 
	.A(FE_OFN1267_router_addr_calc_fft_read_calc_count_9_));
   ADDHXLTS \add_x_22_0/U1_1_8  (.S(\router/addr_calc/fft_read_calc/counter/N54 ), 
	.CO(\add_x_22_0/carry[9] ), 
	.B(\add_x_22_0/carry[8] ), 
	.A(n7571));
   ADDHXLTS \add_x_22_0/U1_1_7  (.S(\router/addr_calc/fft_read_calc/counter/N53 ), 
	.CO(\add_x_22_0/carry[8] ), 
	.B(\add_x_22_0/carry[7] ), 
	.A(n7576));
   ADDHXLTS \add_x_22_0/U1_1_6  (.S(\router/addr_calc/fft_read_calc/counter/N52 ), 
	.CO(\add_x_22_0/carry[7] ), 
	.B(\add_x_22_0/carry[6] ), 
	.A(n7581));
   ADDHXLTS \add_x_22_0/U1_1_5  (.S(\router/addr_calc/fft_read_calc/counter/N51 ), 
	.CO(\add_x_22_0/carry[6] ), 
	.B(\add_x_22_0/carry[5] ), 
	.A(FE_OFN1273_router_addr_calc_fft_read_calc_count_5_));
   ADDHXLTS \add_x_22_0/U1_1_4  (.S(\router/addr_calc/fft_read_calc/counter/N50 ), 
	.CO(\add_x_22_0/carry[5] ), 
	.B(\add_x_22_0/carry[4] ), 
	.A(n7586));
   ADDHXLTS \add_x_22_0/U1_1_3  (.S(\router/addr_calc/fft_read_calc/counter/N49 ), 
	.CO(\add_x_22_0/carry[4] ), 
	.B(\add_x_22_0/carry[3] ), 
	.A(n7591));
   ADDHXLTS \add_x_22_0/U1_1_2  (.S(\router/addr_calc/fft_read_calc/counter/N48 ), 
	.CO(\add_x_22_0/carry[3] ), 
	.B(\add_x_22_0/carry[2] ), 
	.A(n7596));
   INVX2TS U3590 (.Y(n3482), 
	.A(to_fft_empty));
   INVX2TS U3446 (.Y(n3471), 
	.A(to_fir_empty));
   CLKINVX2TS U2649 (.Y(n3769), 
	.A(\fifo_from_fir/tok_xnor_put ));
   INVX2TS U607 (.Y(n3707), 
	.A(\router/ram_write_enable_reg ));
   INVX1TS U951 (.Y(n4004), 
	.A(\fifo_to_fft/tok_xnor_put ));
   CLKINVX1TS U3473 (.Y(n4009), 
	.A(\fifo_to_fft/hang[14] ));
   INVX1TS U2751 (.Y(n3717), 
	.A(\router/iir_write_done ));
   INVX2TS U1433 (.Y(n4025), 
	.A(\router/fir_write_done ));
   INVX1TS U1095 (.Y(n4179), 
	.A(\fifo_to_fir/tok_xnor_put ));
   CLKINVX1TS U3330 (.Y(n4184), 
	.A(\fifo_to_fir/hang[14] ));
   CLKINVX2TS U2018 (.Y(n3789), 
	.A(\fifo_from_fft/tok_xnor_put ));
   INVX2TS U2750 (.Y(\router/addr_calc/iir_write_calc/counter/N212 ), 
	.A(\router/addr_calc/iir_write_calc/counter/hold ));
   CLKINVX2TS U3318 (.Y(n4445), 
	.A(\mips/mips/a/count[0] ));
   NAND4XLTS U602 (.Y(n3704), 
	.D(FE_OFN1273_router_addr_calc_fft_read_calc_count_5_), 
	.C(n7586), 
	.B(n7592), 
	.A(n7487));
   INVX2TS U3872 (.Y(n3850), 
	.A(FE_OFN1283_router_fft_write_done));
   NAND4XLTS U600 (.Y(n3697), 
	.D(FE_OFN1263_router_addr_calc_fft_read_calc_count_16_), 
	.C(n7542), 
	.B(n7547), 
	.A(n7552));
   NAND4XLTS U603 (.Y(n3703), 
	.D(FE_OFN1267_router_addr_calc_fft_read_calc_count_9_), 
	.C(n7572), 
	.B(n7577), 
	.A(n7582));
   NAND4XLTS U373 (.Y(n3567), 
	.D(FE_OFN1248_router_addr_calc_fir_write_calc_count_23_), 
	.C(n7154), 
	.B(n7160), 
	.A(n7166));
   NAND4XLTS U374 (.Y(n3566), 
	.D(n7202), 
	.C(n7206), 
	.B(n7210), 
	.A(FE_OFN1445_router_addr_calc_fir_write_calc_count_0_));
   NAND4XLTS U375 (.Y(n3565), 
	.D(FE_OFN1264_router_addr_calc_fir_write_calc_count_16_), 
	.C(n7184), 
	.B(n7190), 
	.A(n7196));
   NAND4XLTS U377 (.Y(n3572), 
	.D(FE_OFN1272_router_addr_calc_fir_write_calc_count_5_), 
	.C(n7229), 
	.B(n7235), 
	.A(n7118));
   NAND4XLTS U378 (.Y(n3571), 
	.D(\router/addr_calc/fir_write_calc/count[9] ), 
	.C(n7215), 
	.B(n7220), 
	.A(n7225));
   NAND4XLTS U379 (.Y(n3570), 
	.D(FE_OFN1240_router_addr_calc_fir_write_calc_count_27_), 
	.C(n7135), 
	.B(n7142), 
	.A(n7148));
   NAND4XLTS U380 (.Y(n3569), 
	.D(FE_OFN1231_router_addr_calc_fir_write_calc_count_30_), 
	.C(n7240), 
	.B(n7124), 
	.A(n7129));
   NAND4XLTS U604 (.Y(n3702), 
	.D(FE_OFN1237_router_addr_calc_fft_read_calc_count_27_), 
	.C(n7501), 
	.B(n7507), 
	.A(n7512));
   NAND4XLTS U605 (.Y(n3701), 
	.D(FE_OFN1229_router_addr_calc_fft_read_calc_count_30_), 
	.C(n7597), 
	.B(FE_OFN1234_n7492), 
	.A(n7496));
   NAND4XLTS U372 (.Y(n3568), 
	.D(n7244), 
	.C(FE_OFN1261_router_addr_calc_fir_write_calc_count_19_), 
	.B(n7171), 
	.A(n7178));
   NAND4XLTS U529 (.Y(n3658), 
	.D(FE_OFN1238_router_addr_calc_fft_write_calc_count_27_), 
	.C(n7377), 
	.B(n7383), 
	.A(n7388));
   NAND4XLTS U597 (.Y(n3700), 
	.D(n7601), 
	.C(FE_OFN1258_router_addr_calc_fft_read_calc_count_19_), 
	.B(n7531), 
	.A(n7537));
   NAND4XLTS U302 (.Y(n3528), 
	.D(FE_OFN1281_router_addr_calc_iir_write_calc_count_5_), 
	.C(n7095), 
	.B(n7102), 
	.A(n7198));
   NAND4XLTS U303 (.Y(n3527), 
	.D(FE_OFN1280_router_addr_calc_iir_write_calc_count_9_), 
	.C(n7099), 
	.B(n7093), 
	.A(n7090));
   NAND4XLTS U523 (.Y(n3655), 
	.D(FE_OFN1246_router_addr_calc_fft_write_calc_count_23_), 
	.C(n7393), 
	.B(n7398), 
	.A(n7403));
   NAND4XLTS U525 (.Y(n3653), 
	.D(n7418), 
	.C(FE_OFN1270_router_addr_calc_fft_write_calc_count_15_), 
	.B(n7423), 
	.A(n7428));
   NAND4XLTS U304 (.Y(n3526), 
	.D(FE_OFN1439_router_addr_calc_iir_write_calc_count_27_), 
	.C(n7180), 
	.B(n7175), 
	.A(n7169));
   NAND4XLTS U305 (.Y(n3525), 
	.D(\router/addr_calc/iir_write_calc/count[30] ), 
	.C(FE_OFN1825_n7107), 
	.B(n7192), 
	.A(n7186));
   NAND4XLTS U449 (.Y(n3610), 
	.D(n7319), 
	.C(n7324), 
	.B(n7329), 
	.A(\router/addr_calc/fir_read_calc/count[0] ));
   NAND4XLTS U448 (.Y(n3611), 
	.D(FE_OFN1247_router_addr_calc_fir_read_calc_count_23_), 
	.C(n7279), 
	.B(n7284), 
	.A(n7289));
   NAND4XLTS U450 (.Y(n3609), 
	.D(n7304), 
	.C(FE_OFN1271_router_addr_calc_fir_read_calc_count_15_), 
	.B(n7309), 
	.A(n7314));
   NAND4XLTS U452 (.Y(n3616), 
	.D(FE_OFN1276_router_addr_calc_fir_read_calc_count_5_), 
	.C(n7348), 
	.B(n7354), 
	.A(n7249));
   NAND4XLTS U297 (.Y(n3524), 
	.D(n7112), 
	.C(FE_OFN1440_router_addr_calc_iir_write_calc_count_19_), 
	.B(n7144), 
	.A(n7139));
   NAND4XLTS U447 (.Y(n3612), 
	.D(n7363), 
	.C(FE_OFN1260_router_addr_calc_fir_read_calc_count_19_), 
	.B(n7293), 
	.A(n7299));
   NAND4XLTS U453 (.Y(n3615), 
	.D(FE_OFN1269_router_addr_calc_fir_read_calc_count_9_), 
	.C(n7334), 
	.B(n7339), 
	.A(n7344));
   NAND4XLTS U530 (.Y(n3657), 
	.D(FE_OFN1232_n7368), 
	.C(n7478), 
	.B(FE_OFN1233_router_addr_calc_fft_write_calc_count_29_), 
	.A(n7372));
   NAND4XLTS U298 (.Y(n3523), 
	.D(\router/addr_calc/iir_write_calc/count[23] ), 
	.C(n7163), 
	.B(n7157), 
	.A(n7151));
   NAND4XLTS U454 (.Y(n3614), 
	.D(\router/addr_calc/fir_read_calc/count[27] ), 
	.C(n7263), 
	.B(n7269), 
	.A(n7274));
   NAND4XLTS U299 (.Y(n3522), 
	.D(n7116), 
	.C(n7110), 
	.B(n7105), 
	.A(FE_OFN1442_router_addr_calc_iir_write_calc_count_0_));
   NAND4XLTS U455 (.Y(n3613), 
	.D(FE_OFN1230_router_addr_calc_fir_read_calc_count_30_), 
	.C(n7359), 
	.B(FE_OFN1235_n7254), 
	.A(n7258));
   NAND4XLTS U522 (.Y(n3656), 
	.D(n7482), 
	.C(FE_OFN1259_router_addr_calc_fft_write_calc_count_19_), 
	.B(n7407), 
	.A(n7413));
   NAND4XLTS U300 (.Y(n3521), 
	.D(FE_OFN1441_router_addr_calc_iir_write_calc_count_16_), 
	.C(n7133), 
	.B(n7127), 
	.A(n7122));
   NAND4XLTS U599 (.Y(n3698), 
	.D(n7557), 
	.C(n7562), 
	.B(n7567), 
	.A(FE_OFN1444_router_addr_calc_fft_read_calc_count_0_));
   NAND4XLTS U527 (.Y(n3660), 
	.D(n7462), 
	.C(n7467), 
	.B(n7473), 
	.A(FE_OFN1228_router_addr_calc_fft_write_calc_count_31_));
   NAND4XLTS U524 (.Y(n3654), 
	.D(n7433), 
	.C(n7438), 
	.B(n7443), 
	.A(FE_OFN1443_router_addr_calc_fft_write_calc_count_0_));
   NAND4XLTS U528 (.Y(n3659), 
	.D(\router/addr_calc/fft_write_calc/count[9] ), 
	.C(n7448), 
	.B(n7453), 
	.A(n7458));
   NAND4XLTS U598 (.Y(n3699), 
	.D(FE_OFN1245_router_addr_calc_fft_read_calc_count_23_), 
	.C(n7517), 
	.B(n7522), 
	.A(n7527));
   NAND3XLTS U2728 (.Y(n4832), 
	.C(n7603), 
	.B(\router/iir_get_req_reg ), 
	.A(n4830));
   NOR3X1TS U3538 (.Y(n3714), 
	.C(FE_OFN974_n9462), 
	.B(\router/fft_read_done ), 
	.A(\router/fft_write_done ));
   NOR2XLTS U614 (.Y(n3708), 
	.B(n7212), 
	.A(FE_OFN988_n9431));
   AND2XLTS U2713 (.Y(n3472), 
	.B(n9407), 
	.A(FE_OFN978_n9462));
   NAND4BXLTS U613 (.Y(n3716), 
	.D(n3717), 
	.C(n3710), 
	.B(FE_OFN1286_iir_enable), 
	.AN(n3708));
   OAI211X2TS U3871 (.Y(n5346), 
	.C0(\router/fft_get_req_reg ), 
	.B0(n9433), 
	.A1(n3850), 
	.A0(\router/fft_read_done ));
   NAND2XLTS U828 (.Y(n3894), 
	.B(n9498), 
	.A(\fifo_to_fft/fifo_cell13/controller/f_i_put ));
   NAND2XLTS U818 (.Y(n3884), 
	.B(n9498), 
	.A(\fifo_to_fft/fifo_cell15/controller/f_i_put ));
   NAND2XLTS U833 (.Y(n3899), 
	.B(n9498), 
	.A(\fifo_to_fft/fifo_cell12/controller/f_i_put ));
   NAND2XLTS U838 (.Y(n3904), 
	.B(n9499), 
	.A(\fifo_to_fft/fifo_cell11/controller/f_i_put ));
   NAND2XLTS U843 (.Y(n3909), 
	.B(n9497), 
	.A(\fifo_to_fft/fifo_cell10/controller/f_i_put ));
   NAND2XLTS U848 (.Y(n3914), 
	.B(n9499), 
	.A(\fifo_to_fft/fifo_cell9/controller/f_i_put ));
   NAND2XLTS U853 (.Y(n3919), 
	.B(n9499), 
	.A(\fifo_to_fft/fifo_cell8/controller/f_i_put ));
   NAND2XLTS U863 (.Y(n3929), 
	.B(n9499), 
	.A(\fifo_to_fft/fifo_cell6/controller/f_i_put ));
   NAND2XLTS U823 (.Y(n3889), 
	.B(n9498), 
	.A(\fifo_to_fft/fifo_cell14/controller/f_i_put ));
   NAND2XLTS U1628 (.Y(n4517), 
	.B(n9507), 
	.A(\fifo_from_fft/fifo_cell11/controller/f_i_put ));
   NAND2XLTS U1517 (.Y(n4499), 
	.B(n9506), 
	.A(\fifo_from_fft/fifo_cell14/controller/f_i_put ));
   NAND2XLTS U1554 (.Y(n4505), 
	.B(n9507), 
	.A(\fifo_from_fft/fifo_cell13/controller/f_i_put ));
   NAND2XLTS U1665 (.Y(n4523), 
	.B(n9504), 
	.A(\fifo_from_fft/fifo_cell10/controller/f_i_put ));
   NAND2XLTS U1480 (.Y(n4493), 
	.B(n9506), 
	.A(\fifo_from_fft/fifo_cell15/controller/f_i_put ));
   NAND2XLTS U1591 (.Y(n4511), 
	.B(n9506), 
	.A(\fifo_from_fft/fifo_cell12/controller/f_i_put ));
   NAND2XLTS U858 (.Y(n3924), 
	.B(n9500), 
	.A(\fifo_to_fft/fifo_cell7/controller/f_i_put ));
   NAND2XLTS U2185 (.Y(n4691), 
	.B(n9505), 
	.A(\fifo_from_fir/fifo_cell13/controller/f_i_put ));
   NAND2XLTS U962 (.Y(n4059), 
	.B(n9502), 
	.A(\fifo_to_fir/fifo_cell15/controller/f_i_put ));
   NAND2X1TS U967 (.Y(n4064), 
	.B(n9502), 
	.A(\fifo_to_fir/fifo_cell14/controller/f_i_put ));
   NAND2XLTS U972 (.Y(n4069), 
	.B(n9502), 
	.A(\fifo_to_fir/fifo_cell13/controller/f_i_put ));
   NAND2XLTS U977 (.Y(n4074), 
	.B(n9502), 
	.A(\fifo_to_fir/fifo_cell12/controller/f_i_put ));
   NAND2XLTS U868 (.Y(n3934), 
	.B(n9500), 
	.A(\fifo_to_fft/fifo_cell5/controller/f_i_put ));
   NAND2XLTS U982 (.Y(n4079), 
	.B(n9503), 
	.A(\fifo_to_fir/fifo_cell11/controller/f_i_put ));
   NAND2XLTS U987 (.Y(n4084), 
	.B(n9501), 
	.A(\fifo_to_fir/fifo_cell10/controller/f_i_put ));
   NAND2XLTS U873 (.Y(n3939), 
	.B(n9500), 
	.A(\fifo_to_fft/fifo_cell4/controller/f_i_put ));
   NOR2X1TS U1428 (.Y(n4205), 
	.B(acc_done), 
	.A(FE_OFN843_n7619));
   NAND2XLTS U992 (.Y(n4089), 
	.B(n9503), 
	.A(\fifo_to_fir/fifo_cell9/controller/f_i_put ));
   NAND2XLTS U997 (.Y(n4094), 
	.B(n9503), 
	.A(\fifo_to_fir/fifo_cell8/controller/f_i_put ));
   NAND2XLTS U1002 (.Y(n4099), 
	.B(n9504), 
	.A(\fifo_to_fir/fifo_cell7/controller/f_i_put ));
   NAND2XLTS U878 (.Y(n3944), 
	.B(n9501), 
	.A(\fifo_to_fft/fifo_cell3/controller/f_i_put ));
   NAND2XLTS U1007 (.Y(n4104), 
	.B(n9503), 
	.A(\fifo_to_fir/fifo_cell6/controller/f_i_put ));
   NAND2XLTS U883 (.Y(n3949), 
	.B(n9501), 
	.A(\fifo_to_fft/fifo_cell2/controller/f_i_put ));
   NAND2XLTS U1012 (.Y(n4109), 
	.B(n9505), 
	.A(\fifo_to_fir/fifo_cell5/controller/f_i_put ));
   NAND2XLTS U1017 (.Y(n4114), 
	.B(n9504), 
	.A(\fifo_to_fir/fifo_cell4/controller/f_i_put ));
   NAND2XLTS U1022 (.Y(n4119), 
	.B(n9505), 
	.A(\fifo_to_fir/fifo_cell3/controller/f_i_put ));
   NAND2XLTS U888 (.Y(n3954), 
	.B(n9501), 
	.A(\fifo_to_fft/fifo_cell1/controller/f_i_put ));
   NAND2XLTS U895 (.Y(n3960), 
	.B(n9500), 
	.A(\fifo_to_fft/fifo_cell0/controller/f_i_put ));
   NAND2XLTS U1027 (.Y(n4124), 
	.B(n9505), 
	.A(\fifo_to_fir/fifo_cell2/controller/f_i_put ));
   NAND2XLTS U1032 (.Y(n4129), 
	.B(n9506), 
	.A(\fifo_to_fir/fifo_cell1/controller/f_i_put ));
   NAND2XLTS U1039 (.Y(n4135), 
	.B(n9504), 
	.A(\fifo_to_fir/fifo_cell0/controller/f_i_put ));
   NAND2XLTS U1813 (.Y(n4547), 
	.B(n9507), 
	.A(\fifo_from_fft/fifo_cell6/controller/f_i_put ));
   NAND2XLTS U1739 (.Y(n4535), 
	.B(n9507), 
	.A(\fifo_from_fft/fifo_cell8/controller/f_i_put ));
   NOR2X1TS U3322 (.Y(n4444), 
	.B(FE_OFN843_n7619), 
	.A(n4311));
   CLKINVX2TS U1437 (.Y(n4455), 
	.A(n3846));
   INVX1TS U1438 (.Y(n4203), 
	.A(n4456));
   NAND2XLTS U1961 (.Y(n4571), 
	.B(n9508), 
	.A(\fifo_from_fft/fifo_cell2/controller/f_i_put ));
   NAND2XLTS U1776 (.Y(n4541), 
	.B(n9509), 
	.A(\fifo_from_fft/fifo_cell7/controller/f_i_put ));
   NAND2XLTS U2653 (.Y(n4765), 
	.B(n9511), 
	.A(\fifo_from_fir/fifo_cell0/controller/f_i_put ));
   NAND2XLTS U1998 (.Y(n4577), 
	.B(n9510), 
	.A(\fifo_from_fft/fifo_cell1/controller/f_i_put ));
   NAND2XLTS U1887 (.Y(n4559), 
	.B(n9508), 
	.A(\fifo_from_fft/fifo_cell4/controller/f_i_put ));
   NAND2XLTS U2111 (.Y(n4679), 
	.B(n9511), 
	.A(\fifo_from_fir/fifo_cell15/controller/f_i_put ));
   NAND3X1TS U3445 (.Y(n5191), 
	.C(n3471), 
	.B(n9514), 
	.A(FE_OFN1450_acc_fir_get));
   NAND2XLTS U2629 (.Y(n4763), 
	.B(n9513), 
	.A(\fifo_from_fir/fifo_cell1/controller/f_i_put ));
   NAND2XLTS U1924 (.Y(n4565), 
	.B(n9510), 
	.A(\fifo_from_fft/fifo_cell3/controller/f_i_put ));
   NAND3X2TS U3589 (.Y(n5233), 
	.C(n3482), 
	.B(n9514), 
	.A(FE_OFN1448_acc_fft_get));
   NAND2XLTS U2022 (.Y(n4579), 
	.B(n9508), 
	.A(\fifo_from_fft/fifo_cell0/controller/f_i_put ));
   NAND2XLTS U1850 (.Y(n4553), 
	.B(n9509), 
	.A(\fifo_from_fft/fifo_cell5/controller/f_i_put ));
   NAND2XLTS U2259 (.Y(n4703), 
	.B(n9512), 
	.A(\fifo_from_fir/fifo_cell11/controller/f_i_put ));
   NAND2XLTS U2407 (.Y(n4727), 
	.B(n9512), 
	.A(\fifo_from_fir/fifo_cell7/controller/f_i_put ));
   NAND2XLTS U2370 (.Y(n4721), 
	.B(n9511), 
	.A(\fifo_from_fir/fifo_cell8/controller/f_i_put ));
   NAND2XLTS U2444 (.Y(n4733), 
	.B(n9510), 
	.A(\fifo_from_fir/fifo_cell6/controller/f_i_put ));
   NAND2XLTS U2296 (.Y(n4709), 
	.B(n9509), 
	.A(\fifo_from_fir/fifo_cell10/controller/f_i_put ));
   NAND2XLTS U2222 (.Y(n4697), 
	.B(n9510), 
	.A(\fifo_from_fir/fifo_cell12/controller/f_i_put ));
   NAND2XLTS U2481 (.Y(n4739), 
	.B(n9513), 
	.A(\fifo_from_fir/fifo_cell5/controller/f_i_put ));
   NAND2XLTS U2518 (.Y(n4745), 
	.B(n9511), 
	.A(\fifo_from_fir/fifo_cell4/controller/f_i_put ));
   NAND2XLTS U2592 (.Y(n4757), 
	.B(n9512), 
	.A(\fifo_from_fir/fifo_cell2/controller/f_i_put ));
   NOR3X1TS U3870 (.Y(n4643), 
	.C(n5346), 
	.B(from_fft_empty), 
	.A(FE_OFN795_n7619));
   NAND2XLTS U2148 (.Y(n4685), 
	.B(n9509), 
	.A(\fifo_from_fir/fifo_cell14/controller/f_i_put ));
   NAND2XLTS U2555 (.Y(n4751), 
	.B(n9513), 
	.A(\fifo_from_fir/fifo_cell3/controller/f_i_put ));
   NAND2XLTS U1702 (.Y(n4529), 
	.B(n9508), 
	.A(\fifo_from_fft/fifo_cell9/controller/f_i_put ));
   NAND2XLTS U2333 (.Y(n4715), 
	.B(n9512), 
	.A(\fifo_from_fir/fifo_cell9/controller/f_i_put ));
   AOI21X1TS U606 (.Y(FE_OFN848_ram_write_enable), 
	.B0(n3707), 
	.A1(n3706), 
	.A0(n3705));
   NAND3XLTS U1432 (.Y(n4454), 
	.C(n4455), 
	.B(n7960), 
	.A(FE_OFN1283_router_fft_write_done));
   NOR3BXLTS U3474 (.Y(\fifo_to_fft/fifo_cell15/N7 ), 
	.C(n5233), 
	.B(\fifo_to_fft/fifo_cell15/control_signal ), 
	.AN(\fifo_to_fft/fifo_cell15/reg_gtok/token ));
   CLKINVX2TS U3444 (.Y(n4134), 
	.A(n5191));
   INVX2TS U3588 (.Y(n3959), 
	.A(n5233));
   NOR3BXLTS U3331 (.Y(\fifo_to_fir/fifo_cell15/N7 ), 
	.C(n5191), 
	.B(\fifo_to_fir/fifo_cell15/control_signal ), 
	.AN(\fifo_to_fir/fifo_cell15/reg_gtok/token ));
   NOR3X1TS U3815 (.Y(n5326), 
	.C(\fifo_from_fft/fifo_cell1/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell1/controller/write_enable ), 
	.A(n7524));
   OAI31XLTS U1431 (.Y(n4453), 
	.B0(n4454), 
	.A2(n4200), 
	.A1(n7212), 
	.A0(n4025));
   NAND2XLTS U1104 (.Y(n4201), 
	.B(n3846), 
	.A(n4202));
   NAND4BXLTS U810 (.Y(n3847), 
	.D(n3849), 
	.C(n9480), 
	.B(n9434), 
	.AN(n3848));
   NOR2XLTS U227 (.Y(n3480), 
	.B(n7607), 
	.A(n3472));
   NAND2XLTS U217 (.Y(n3463), 
	.B(n3467), 
	.A(n7203));
   NAND2XLTS U1422 (.Y(n4442), 
	.B(\mips/mips/a/countflag ), 
	.A(\mips/mips/a/count[0] ));
   NAND2X1TS U3726 (.Y(n4764), 
	.B(\fifo_from_fir/fifo_cell0/reg_gtok/token ), 
	.A(FE_OFN735_n4829));
   NOR3X1TS U3782 (.Y(n5318), 
	.C(\fifo_from_fft/fifo_cell9/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell9/controller/write_enable ), 
	.A(n7485));
   NOR3X1TS U3766 (.Y(n5314), 
	.C(\fifo_from_fft/fifo_cell13/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell13/controller/write_enable ), 
	.A(n7465));
   NOR3X1TS U3774 (.Y(n5316), 
	.C(\fifo_from_fft/fifo_cell11/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell11/controller/write_enable ), 
	.A(n7475));
   NOR3X1TS U3762 (.Y(n5313), 
	.C(\fifo_from_fft/fifo_cell14/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell14/controller/write_enable ), 
	.A(n7460));
   NOR3X1TS U3770 (.Y(n5315), 
	.C(\fifo_from_fft/fifo_cell12/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell12/controller/write_enable ), 
	.A(n7470));
   NAND2XLTS U3837 (.Y(n4500), 
	.B(\fifo_from_fft/fifo_cell13/reg_gtok/token ), 
	.A(FE_OFN723_n4643));
   NAND2XLTS U3843 (.Y(n4494), 
	.B(\fifo_from_fft/fifo_cell14/reg_gtok/token ), 
	.A(FE_OFN725_n4643));
   NOR3X1TS U3794 (.Y(n5321), 
	.C(\fifo_from_fft/fifo_cell6/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell6/controller/write_enable ), 
	.A(n7499));
   NOR3X1TS U3639 (.Y(n5279), 
	.C(\fifo_from_fir/fifo_cell9/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell9/controller/write_enable ), 
	.A(n7559));
   NOR3X1TS U3635 (.Y(n5278), 
	.C(\fifo_from_fir/fifo_cell10/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell10/controller/write_enable ), 
	.A(n7554));
   NOR3X1TS U3651 (.Y(n5282), 
	.C(\fifo_from_fir/fifo_cell6/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell6/controller/write_enable ), 
	.A(n7574));
   NOR3X1TS U3790 (.Y(n5320), 
	.C(\fifo_from_fft/fifo_cell7/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell7/controller/write_enable ), 
	.A(n7494));
   NOR3X1TS U3619 (.Y(n5274), 
	.C(\fifo_from_fir/fifo_cell14/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell14/controller/write_enable ), 
	.A(n7534));
   NOR3X1TS U3647 (.Y(n5281), 
	.C(\fifo_from_fir/fifo_cell7/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell7/controller/write_enable ), 
	.A(n7569));
   NOR3X1TS U3802 (.Y(n5323), 
	.C(\fifo_from_fft/fifo_cell4/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell4/controller/write_enable ), 
	.A(n7509));
   NOR3X1TS U3623 (.Y(n5275), 
	.C(\fifo_from_fir/fifo_cell13/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell13/controller/write_enable ), 
	.A(n7539));
   NOR3X1TS U3627 (.Y(n5276), 
	.C(\fifo_from_fir/fifo_cell12/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell12/controller/write_enable ), 
	.A(n7544));
   NOR3X1TS U3655 (.Y(n5283), 
	.C(\fifo_from_fir/fifo_cell5/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell5/controller/write_enable ), 
	.A(n7579));
   NOR3X1TS U3659 (.Y(n5284), 
	.C(\fifo_from_fir/fifo_cell4/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell4/controller/write_enable ), 
	.A(n7584));
   NOR3X1TS U3663 (.Y(n5285), 
	.C(\fifo_from_fir/fifo_cell3/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell3/controller/write_enable ), 
	.A(n7589));
   NOR3X1TS U3806 (.Y(n5324), 
	.C(\fifo_from_fft/fifo_cell3/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell3/controller/write_enable ), 
	.A(n7514));
   NOR3X1TS U3798 (.Y(n5322), 
	.C(\fifo_from_fft/fifo_cell5/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell5/controller/write_enable ), 
	.A(n7504));
   NOR3X1TS U3672 (.Y(n5287), 
	.C(\fifo_from_fir/fifo_cell1/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell1/controller/write_enable ), 
	.A(n7599));
   NOR3X1TS U3631 (.Y(n5277), 
	.C(\fifo_from_fir/fifo_cell11/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell11/controller/write_enable ), 
	.A(n7549));
   NOR3X1TS U3778 (.Y(n5317), 
	.C(\fifo_from_fft/fifo_cell10/controller/valid_read ), 
	.B(\fifo_from_fft/fifo_cell10/controller/write_enable ), 
	.A(n7480));
   NOR3X1TS U3667 (.Y(n5286), 
	.C(\fifo_from_fir/fifo_cell2/controller/valid_read ), 
	.B(\fifo_from_fir/fifo_cell2/controller/write_enable ), 
	.A(n7594));
   NAND2XLTS U3694 (.Y(n4686), 
	.B(\fifo_from_fir/fifo_cell13/reg_gtok/token ), 
	.A(FE_OFN742_n4829));
   NAND2X1TS U3700 (.Y(n4680), 
	.B(\fifo_from_fir/fifo_cell14/reg_gtok/token ), 
	.A(FE_OFN742_n4829));
   OAI2BB1XLTS U2693 (.Y(n6754), 
	.B0(n4734), 
	.A1N(n7966), 
	.A0N(\fifo_from_fir/fifo_cell6/reg_gtok/token ));
   OAI2BB1XLTS U2694 (.Y(n6755), 
	.B0(n4740), 
	.A1N(n7966), 
	.A0N(\fifo_from_fir/fifo_cell5/reg_gtok/token ));
   OAI2BB1XLTS U2695 (.Y(n6756), 
	.B0(n4746), 
	.A1N(n7965), 
	.A0N(\fifo_from_fir/fifo_cell4/reg_gtok/token ));
   OAI2BB1XLTS U2698 (.Y(n6759), 
	.B0(n4764), 
	.A1N(n7963), 
	.A0N(\fifo_from_fir/fifo_cell1/reg_gtok/token ));
   OAI2BB1XLTS U2061 (.Y(n6224), 
	.B0(n4542), 
	.A1N(n7970), 
	.A0N(\fifo_from_fft/fifo_cell7/reg_gtok/token ));
   OAI2BB1XLTS U2063 (.Y(n6226), 
	.B0(n4554), 
	.A1N(n7971), 
	.A0N(\fifo_from_fft/fifo_cell5/reg_gtok/token ));
   OAI2BB1XLTS U2064 (.Y(n6227), 
	.B0(n4560), 
	.A1N(n7969), 
	.A0N(\fifo_from_fft/fifo_cell4/reg_gtok/token ));
   OAI2BB1XLTS U2060 (.Y(n6223), 
	.B0(n4536), 
	.A1N(n7971), 
	.A0N(\fifo_from_fft/fifo_cell8/reg_gtok/token ));
   OAI2BB1XLTS U2065 (.Y(n6228), 
	.B0(n4566), 
	.A1N(n7968), 
	.A0N(\fifo_from_fft/fifo_cell3/reg_gtok/token ));
   OAI2BB1XLTS U2066 (.Y(n6229), 
	.B0(n4572), 
	.A1N(n7971), 
	.A0N(\fifo_from_fft/fifo_cell2/reg_gtok/token ));
   OAI2BB1XLTS U2059 (.Y(n6222), 
	.B0(n4530), 
	.A1N(n7969), 
	.A0N(\fifo_from_fft/fifo_cell9/reg_gtok/token ));
   OAI2BB1XLTS U2067 (.Y(n6230), 
	.B0(n4578), 
	.A1N(n7968), 
	.A0N(\fifo_from_fft/fifo_cell1/reg_gtok/token ));
   OAI2BB1XLTS U2058 (.Y(n6221), 
	.B0(n4524), 
	.A1N(n7970), 
	.A0N(\fifo_from_fft/fifo_cell10/reg_gtok/token ));
   OAI2BB1XLTS U2057 (.Y(n6220), 
	.B0(n4518), 
	.A1N(n7971), 
	.A0N(\fifo_from_fft/fifo_cell11/reg_gtok/token ));
   OAI2BB1XLTS U2056 (.Y(n6219), 
	.B0(n4512), 
	.A1N(n7968), 
	.A0N(\fifo_from_fft/fifo_cell12/reg_gtok/token ));
   OAI2BB1XLTS U2054 (.Y(n6217), 
	.B0(n4500), 
	.A1N(n7970), 
	.A0N(\fifo_from_fft/fifo_cell14/reg_gtok/token ));
   OAI2BB1XLTS U2053 (.Y(n6216), 
	.B0(n4494), 
	.A1N(n7970), 
	.A0N(\fifo_from_fft/fifo_cell15/reg_gtok/token ));
   OAI2BB1XLTS U2055 (.Y(n6218), 
	.B0(n4506), 
	.A1N(n7969), 
	.A0N(\fifo_from_fft/fifo_cell13/reg_gtok/token ));
   OAI2BB1XLTS U2062 (.Y(n6225), 
	.B0(n4548), 
	.A1N(n7969), 
	.A0N(\fifo_from_fft/fifo_cell6/reg_gtok/token ));
   OAI2BB1XLTS U2697 (.Y(n6758), 
	.B0(n4758), 
	.A1N(n7964), 
	.A0N(\fifo_from_fir/fifo_cell2/reg_gtok/token ));
   OAI2BB1XLTS U2696 (.Y(n6757), 
	.B0(n4752), 
	.A1N(n7964), 
	.A0N(\fifo_from_fir/fifo_cell3/reg_gtok/token ));
   OAI2BB1XLTS U2692 (.Y(n6753), 
	.B0(n4728), 
	.A1N(n7965), 
	.A0N(\fifo_from_fir/fifo_cell7/reg_gtok/token ));
   AOI21X1TS U1420 (.Y(n5700), 
	.B0(n4443), 
	.A1(n4442), 
	.A0(n4441));
   OAI2BB1XLTS U2691 (.Y(n6752), 
	.B0(n4722), 
	.A1N(n7965), 
	.A0N(\fifo_from_fir/fifo_cell8/reg_gtok/token ));
   OAI2BB1XLTS U2690 (.Y(n6751), 
	.B0(n4716), 
	.A1N(n7964), 
	.A0N(\fifo_from_fir/fifo_cell9/reg_gtok/token ));
   OAI2BB1XLTS U2689 (.Y(n6750), 
	.B0(n4710), 
	.A1N(n7966), 
	.A0N(\fifo_from_fir/fifo_cell10/reg_gtok/token ));
   OAI2BB1XLTS U2688 (.Y(n6749), 
	.B0(n4704), 
	.A1N(n7966), 
	.A0N(\fifo_from_fir/fifo_cell11/reg_gtok/token ));
   OAI2BB1XLTS U2687 (.Y(n6748), 
	.B0(n4698), 
	.A1N(n7963), 
	.A0N(\fifo_from_fir/fifo_cell12/reg_gtok/token ));
   OAI2BB1XLTS U2686 (.Y(n6747), 
	.B0(n4692), 
	.A1N(n7963), 
	.A0N(\fifo_from_fir/fifo_cell13/reg_gtok/token ));
   OAI2BB1XLTS U2685 (.Y(n6746), 
	.B0(n4686), 
	.A1N(n7964), 
	.A0N(\fifo_from_fir/fifo_cell14/reg_gtok/token ));
   OAI2BB1XLTS U2684 (.Y(n6745), 
	.B0(n4680), 
	.A1N(n7965), 
	.A0N(\fifo_from_fir/fifo_cell15/reg_gtok/token ));
   INVX2TS U3323 (.Y(from_fir_full), 
	.A(n3465));
   AOI22XLTS U3414 (.Y(n5219), 
	.B1(n4103), 
	.B0(n4108), 
	.A1(\fifo_to_fir/fifo_cell5/data_out/N35 ), 
	.A0(\fifo_to_fir/fifo_cell6/data_out/N35 ));
   CLKINVX1TS U795 (.Y(n3476), 
	.A(n3484));
   AOI22XLTS U3558 (.Y(n5261), 
	.B1(n3928), 
	.B0(n3933), 
	.A1(\fifo_to_fft/fifo_cell5/data_out/N35 ), 
	.A0(\fifo_to_fft/fifo_cell6/data_out/N35 ));
   NAND2XLTS U2721 (.Y(n3835), 
	.B(n3484), 
	.A(\router/data_cntl/fft_full_flag ));
   NAND2XLTS U230 (.Y(n3483), 
	.B(n3477), 
	.A(n3484));
   AND2XLTS U3434 (.Y(n4058), 
	.B(FE_OFN684_n4134), 
	.A(\fifo_to_fir/fifo_cell14/reg_gtok/token ));
   AND2XLTS U3443 (.Y(n4128), 
	.B(FE_OFN683_n4134), 
	.A(\fifo_to_fir/fifo_cell0/reg_gtok/token ));
   AND2XLTS U3578 (.Y(n3883), 
	.B(n3959), 
	.A(\fifo_to_fft/fifo_cell14/reg_gtok/token ));
   INVX2TS U3324 (.Y(from_fft_full), 
	.A(n3477));
   AND2XLTS U3587 (.Y(n3953), 
	.B(FE_OFN700_n3959), 
	.A(\fifo_to_fft/fifo_cell0/reg_gtok/token ));
   OAI32XLTS U1423 (.Y(n5701), 
	.B1(n8051), 
	.B0(n4445), 
	.A2(\mips/mips/a/N49 ), 
	.A1(\mips/mips/a/count[0] ), 
	.A0(n9370));
   NOR2BXLTS U794 (.Y(n3830), 
	.B(n3835), 
	.AN(n3834));
   AOI32XLTS U226 (.Y(n3481), 
	.B1(n9433), 
	.B0(n3483), 
	.A2(FE_OFN1217_n3478), 
	.A1(n9433), 
	.A0(n3482));
   AOI22XLTS U3409 (.Y(n5220), 
	.B1(n4113), 
	.B0(n4118), 
	.A1(\fifo_to_fir/fifo_cell3/data_out/N35 ), 
	.A0(\fifo_to_fir/fifo_cell4/data_out/N35 ));
   OAI2BB1XLTS U821 (.Y(n5472), 
	.B0(n3888), 
	.A1N(n7974), 
	.A0N(\fifo_to_fft/fifo_cell14/reg_gtok/token ));
   AOI22XLTS U3437 (.Y(n5225), 
	.B1(n4073), 
	.B0(n4078), 
	.A1(\fifo_to_fir/fifo_cell11/data_out/N35 ), 
	.A0(\fifo_to_fir/fifo_cell12/data_out/N35 ));
   INVX1TS U228 (.Y(n3479), 
	.A(\router/data_cntl/N135 ));
   AOI22XLTS U3426 (.Y(n5223), 
	.B1(n4098), 
	.B0(n4063), 
	.A1(\fifo_to_fir/fifo_cell14/data_out/N35 ), 
	.A0(\fifo_to_fir/fifo_cell7/data_out/N35 ));
   CLKINVX1TS U178 (.Y(n2848), 
	.A(n3830));
   AOI22XLTS U3421 (.Y(n5224), 
	.B1(n4088), 
	.B0(n4093), 
	.A1(\fifo_to_fir/fifo_cell8/data_out/N35 ), 
	.A0(\fifo_to_fir/fifo_cell9/data_out/N35 ));
   OAI2BB1XLTS U846 (.Y(n5487), 
	.B0(n3913), 
	.A1N(n7974), 
	.A0N(\fifo_to_fft/fifo_cell9/reg_gtok/token ));
   NAND2XLTS U798 (.Y(n3837), 
	.B(n7608), 
	.A(\router/data_cntl/fir_full_flag ));
   AOI22XLTS U3565 (.Y(n5266), 
	.B1(n3913), 
	.B0(n3918), 
	.A1(\fifo_to_fft/fifo_cell8/data_out/N35 ), 
	.A0(\fifo_to_fft/fifo_cell9/data_out/N35 ));
   OAI2BB1XLTS U841 (.Y(n5484), 
	.B0(n3908), 
	.A1N(n7976), 
	.A0N(\fifo_to_fft/fifo_cell10/reg_gtok/token ));
   NAND2XLTS U222 (.Y(n3473), 
	.B(n3465), 
	.A(n7609));
   OAI2BB1XLTS U881 (.Y(n5508), 
	.B0(n3948), 
	.A1N(n7974), 
	.A0N(\fifo_to_fft/fifo_cell2/reg_gtok/token ));
   OAI2BB1XLTS U831 (.Y(n5478), 
	.B0(n3898), 
	.A1N(n7973), 
	.A0N(\fifo_to_fft/fifo_cell12/reg_gtok/token ));
   OAI2BB1XLTS U826 (.Y(n5475), 
	.B0(n3893), 
	.A1N(n7973), 
	.A0N(\fifo_to_fft/fifo_cell13/reg_gtok/token ));
   OAI2BB1XLTS U851 (.Y(n5490), 
	.B0(n3918), 
	.A1N(n7975), 
	.A0N(\fifo_to_fft/fifo_cell8/reg_gtok/token ));
   AOI22XLTS U3581 (.Y(n5267), 
	.B1(n3898), 
	.B0(n3903), 
	.A1(\fifo_to_fft/fifo_cell11/data_out/N35 ), 
	.A0(\fifo_to_fft/fifo_cell12/data_out/N35 ));
   OAI2BB1XLTS U856 (.Y(n5493), 
	.B0(n3923), 
	.A1N(n7975), 
	.A0N(\fifo_to_fft/fifo_cell7/reg_gtok/token ));
   AOI22XLTS U3570 (.Y(n5265), 
	.B1(n3923), 
	.B0(n3888), 
	.A1(\fifo_to_fft/fifo_cell14/data_out/N35 ), 
	.A0(\fifo_to_fft/fifo_cell7/data_out/N35 ));
   OAI2BB1XLTS U866 (.Y(n5499), 
	.B0(n3933), 
	.A1N(n7976), 
	.A0N(\fifo_to_fft/fifo_cell5/reg_gtok/token ));
   OAI2BB1XLTS U836 (.Y(n5481), 
	.B0(n3903), 
	.A1N(n7976), 
	.A0N(\fifo_to_fft/fifo_cell11/reg_gtok/token ));
   AOI22XLTS U3553 (.Y(n5262), 
	.B1(n3938), 
	.B0(n3943), 
	.A1(\fifo_to_fft/fifo_cell3/data_out/N35 ), 
	.A0(\fifo_to_fft/fifo_cell4/data_out/N35 ));
   OAI2BB1XLTS U876 (.Y(n5505), 
	.B0(n3943), 
	.A1N(n7974), 
	.A0N(\fifo_to_fft/fifo_cell3/reg_gtok/token ));
   OAI2BB1XLTS U871 (.Y(n5502), 
	.B0(n3938), 
	.A1N(n7975), 
	.A0N(\fifo_to_fft/fifo_cell4/reg_gtok/token ));
   OAI2BB1XLTS U861 (.Y(n5496), 
	.B0(n3928), 
	.A1N(n7976), 
	.A0N(\fifo_to_fft/fifo_cell6/reg_gtok/token ));
   OAI2BB1XLTS U1010 (.Y(n5551), 
	.B0(n4108), 
	.A1N(n7615), 
	.A0N(\fifo_to_fir/fifo_cell5/reg_gtok/token ));
   OAI2BB1XLTS U985 (.Y(n5536), 
	.B0(n4083), 
	.A1N(n7614), 
	.A0N(\fifo_to_fir/fifo_cell10/reg_gtok/token ));
   OAI2BB1XLTS U1025 (.Y(n5560), 
	.B0(n4123), 
	.A1N(n7614), 
	.A0N(\fifo_to_fir/fifo_cell2/reg_gtok/token ));
   OAI2BB1XLTS U1005 (.Y(n5548), 
	.B0(n4103), 
	.A1N(n7614), 
	.A0N(\fifo_to_fir/fifo_cell6/reg_gtok/token ));
   OAI2BB1XLTS U886 (.Y(n5511), 
	.B0(n7335), 
	.A1N(n7973), 
	.A0N(\fifo_to_fft/fifo_cell1/reg_gtok/token ));
   OAI2BB1XLTS U1000 (.Y(n5545), 
	.B0(n4098), 
	.A1N(n7617), 
	.A0N(\fifo_to_fir/fifo_cell7/reg_gtok/token ));
   CLKINVX1TS U3577 (.Y(\fifo_to_fft/fifo_cell15/data_out/N35 ), 
	.A(n7236));
   OAI2BB1XLTS U970 (.Y(n5527), 
	.B0(n4068), 
	.A1N(n7615), 
	.A0N(\fifo_to_fir/fifo_cell13/reg_gtok/token ));
   OAI2BB1XLTS U1030 (.Y(n5563), 
	.B0(n7444), 
	.A1N(n7615), 
	.A0N(\fifo_to_fir/fifo_cell1/reg_gtok/token ));
   OAI2BB1XLTS U990 (.Y(n5539), 
	.B0(n4088), 
	.A1N(n7615), 
	.A0N(\fifo_to_fir/fifo_cell9/reg_gtok/token ));
   OAI2BB1XLTS U1020 (.Y(n5557), 
	.B0(n4118), 
	.A1N(n7617), 
	.A0N(\fifo_to_fir/fifo_cell3/reg_gtok/token ));
   OAI2BB1XLTS U995 (.Y(n5542), 
	.B0(n4093), 
	.A1N(n7616), 
	.A0N(\fifo_to_fir/fifo_cell8/reg_gtok/token ));
   OAI2BB1XLTS U1015 (.Y(n5554), 
	.B0(n4113), 
	.A1N(n7616), 
	.A0N(\fifo_to_fir/fifo_cell4/reg_gtok/token ));
   NOR2XLTS U797 (.Y(n3825), 
	.B(n3838), 
	.A(n3837));
   AOI32XLTS U221 (.Y(n3468), 
	.B1(n7203), 
	.B0(n3473), 
	.A2(n3467), 
	.A1(n7203), 
	.A0(n3471));
   OAI2BB1XLTS U965 (.Y(n5524), 
	.B0(n4063), 
	.A1N(n7614), 
	.A0N(\fifo_to_fir/fifo_cell14/reg_gtok/token ));
   OAI2BB1XLTS U980 (.Y(n5533), 
	.B0(n4078), 
	.A1N(n7617), 
	.A0N(\fifo_to_fir/fifo_cell11/reg_gtok/token ));
   OAI2BB1XLTS U975 (.Y(n5530), 
	.B0(n4073), 
	.A1N(n7616), 
	.A0N(\fifo_to_fir/fifo_cell12/reg_gtok/token ));
   OAI2BB1XLTS U960 (.Y(n5521), 
	.B0(n7345), 
	.A1N(n7617), 
	.A0N(\fifo_to_fir/fifo_cell15/reg_gtok/token ));
   CLKINVX1TS U3433 (.Y(\fifo_to_fir/fifo_cell15/data_out/N35 ), 
	.A(n7345));
   OAI2BB1XLTS U816 (.Y(n5469), 
	.B0(n7236), 
	.A1N(n7975), 
	.A0N(\fifo_to_fft/fifo_cell15/reg_gtok/token ));
   NOR2X1TS U2718 (.Y(n3829), 
	.B(n3839), 
	.A(\router/data_cntl/N151 ));
   AOI22XLTS U3576 (.Y(n5268), 
	.B1(n3908), 
	.B0(n7237), 
	.A1(\fifo_to_fft/fifo_cell15/data_out/N35 ), 
	.A0(\fifo_to_fft/fifo_cell10/data_out/N35 ));
   AOI22XLTS U3547 (.Y(n5260), 
	.B1(n7336), 
	.B0(n3893), 
	.A1(\fifo_to_fft/fifo_cell13/data_out/N35 ), 
	.A0(\fifo_to_fft/fifo_cell1/data_out/N35 ));
   AOI22XLTS U3403 (.Y(n5218), 
	.B1(n7445), 
	.B0(n4068), 
	.A1(\fifo_to_fir/fifo_cell13/data_out/N35 ), 
	.A0(\fifo_to_fir/fifo_cell1/data_out/N35 ));
   AOI22XLTS U3432 (.Y(n5226), 
	.B1(n4083), 
	.B0(n7346), 
	.A1(\fifo_to_fir/fifo_cell15/data_out/N35 ), 
	.A0(\fifo_to_fir/fifo_cell10/data_out/N35 ));
   AOI211XLTS U219 (.Y(n3469), 
	.C0(n7606), 
	.B0(n9432), 
	.A1(n3470), 
	.A0(\router/data_cntl/N137 ));
   AOI22X1TS U290 (.Y(n3516), 
	.B1(\router/addr_calc/iir_write_calc/counter/N48 ), 
	.B0(FE_OFN938_n3487), 
	.A1(FE_OFN942_n3486), 
	.A0(FE_OFN1825_n7107));
   AOI22X1TS U294 (.Y(n3518), 
	.B1(n7959), 
	.B0(FE_OFN937_n3487), 
	.A1(FE_OFN945_n3486), 
	.A0(\router/addr_calc/iir_write_calc/count[0] ));
   AOI22X1TS U286 (.Y(n3514), 
	.B1(\router/addr_calc/iir_write_calc/counter/N50 ), 
	.B0(FE_OFN939_n3487), 
	.A1(FE_OFN942_n3486), 
	.A0(n7095));
   AOI22X1TS U280 (.Y(n3511), 
	.B1(\router/addr_calc/iir_write_calc/counter/N53 ), 
	.B0(FE_OFN937_n3487), 
	.A1(FE_OFN947_n3486), 
	.A0(n7092));
   AOI22X1TS U282 (.Y(n3512), 
	.B1(\router/addr_calc/iir_write_calc/counter/N52 ), 
	.B0(FE_OFN937_n3487), 
	.A1(FE_OFN945_n3486), 
	.A0(n7089));
   AOI22X1TS U292 (.Y(n3517), 
	.B1(\router/addr_calc/iir_write_calc/counter/N47 ), 
	.B0(FE_OFN938_n3487), 
	.A1(FE_OFN945_n3486), 
	.A0(n7112));
   AOI22X1TS U266 (.Y(n3504), 
	.B1(\router/addr_calc/iir_write_calc/counter/N60 ), 
	.B0(FE_OFN934_n3487), 
	.A1(FE_OFN949_n3486), 
	.A0(n7126));
   AOI22X1TS U268 (.Y(n3505), 
	.B1(\router/addr_calc/iir_write_calc/counter/N59 ), 
	.B0(FE_OFN935_n3487), 
	.A1(FE_OFN949_n3486), 
	.A0(n7121));
   AOI22X1TS U284 (.Y(n3513), 
	.B1(\router/addr_calc/iir_write_calc/counter/N51 ), 
	.B0(FE_OFN939_n3487), 
	.A1(FE_OFN940_n3486), 
	.A0(FE_OFN1281_router_addr_calc_iir_write_calc_count_5_));
   OAI2BB1XLTS U2068 (.Y(n6231), 
	.B0(n4580), 
	.A1N(n7968), 
	.A0N(\fifo_from_fft/fifo_cell0/reg_gtok/token ));
   AND4XLTS U790 (.Y(n3827), 
	.D(n9391), 
	.C(FE_OFN988_n9431), 
	.B(FE_OFN976_n9462), 
	.A(n3829));
   INVX1TS U3825 (.Y(\fifo_from_fft/fifo_cell0/data_out/N35 ), 
	.A(n4580));
   OAI2BB1XLTS U2699 (.Y(n6760), 
	.B0(n4766), 
	.A1N(n7963), 
	.A0N(\fifo_from_fir/fifo_cell0/reg_gtok/token ));
   NAND2XLTS U273 (.Y(\router/addr_calc/iir_write_calc/counter/N188 ), 
	.B(n3508), 
	.A(FE_OFN1298_iir_enable));
   NOR3X1TS U2071 (.Y(n3758), 
	.C(n3755), 
	.B(n3840), 
	.A(\router/data_to_fft ));
   INVX1TS U3682 (.Y(\fifo_from_fir/fifo_cell0/data_out/N35 ), 
	.A(n4766));
   AOI22X1TS U264 (.Y(n3503), 
	.B1(\router/addr_calc/iir_write_calc/counter/N61 ), 
	.B0(FE_OFN934_n3487), 
	.A1(FE_OFN949_n3486), 
	.A0(n7132));
   NAND2XLTS U271 (.Y(\router/addr_calc/iir_write_calc/counter/N189 ), 
	.B(n3507), 
	.A(FE_OFN1298_iir_enable));
   NAND2XLTS U269 (.Y(\router/addr_calc/iir_write_calc/counter/N190 ), 
	.B(n3506), 
	.A(FE_OFN1294_iir_enable));
   NAND2XLTS U287 (.Y(\router/addr_calc/iir_write_calc/counter/N181 ), 
	.B(n3515), 
	.A(FE_OFN1300_iir_enable));
   NAND2XLTS U277 (.Y(\router/addr_calc/iir_write_calc/counter/N186 ), 
	.B(n3510), 
	.A(FE_OFN1299_iir_enable));
   NAND2XLTS U275 (.Y(\router/addr_calc/iir_write_calc/counter/N187 ), 
	.B(n3509), 
	.A(FE_OFN1298_iir_enable));
   OAI31XLTS U791 (.Y(n3831), 
	.B0(n3832), 
	.A2(n3476), 
	.A1(n7611), 
	.A0(FE_OFN979_n9462));
   AO21XLTS U2704 (.Y(n6762), 
	.B0(n3757), 
	.A1(n4832), 
	.A0(\router/iir_get_req_reg ));
   AO21XLTS U2070 (.Y(n6232), 
	.B0(n3758), 
	.A1(\router/fft_get_req_reg ), 
	.A0(\router/ram_read_enable_reg ));
   AOI22X1TS U262 (.Y(n3502), 
	.B1(\router/addr_calc/iir_write_calc/counter/N62 ), 
	.B0(FE_OFN934_n3487), 
	.A1(FE_OFN950_n3486), 
	.A0(FE_OFN1441_router_addr_calc_iir_write_calc_count_16_));
   OAI21X1TS U2628 (.Y(n4761), 
	.B0(FE_OFN666_n4759), 
	.A1(n4764), 
	.A0(n7599));
   OAI21XLTS U1997 (.Y(n4575), 
	.B0(n4573), 
	.A1(n4578), 
	.A0(n7524));
   NAND2XLTS U808 (.Y(n3845), 
	.B(n3843), 
	.A(\router/data_from_fir ));
   NAND4XLTS U807 (.Y(n3844), 
	.D(FE_OFN978_n9462), 
	.C(\router/data_to_fir ), 
	.B(\router/data_from_fir ), 
	.A(n9406));
   AOI22X1TS U260 (.Y(n3501), 
	.B1(\router/addr_calc/iir_write_calc/counter/N63 ), 
	.B0(FE_OFN932_n3487), 
	.A1(FE_OFN950_n3486), 
	.A0(n7138));
   AO22XLTS U2618 (.Y(n6735), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[6] ), 
	.B0(FE_OFN345_n4760), 
	.A1(FE_OFN1774_acc_fir_data_in_6_), 
	.A0(FE_OFN668_n4759));
   OAI21X1TS U3399 (.Y(n4133), 
	.B0(FE_OFN683_n4134), 
	.A1(n5213), 
	.A0(\fifo_to_fir/fifo_cell15/reg_gtok/token ));
   OAI21XLTS U1996 (.Y(n6214), 
	.B0(n4575), 
	.A1(n4577), 
	.A0(\fifo_from_fft/fifo_cell1/data_out/N35 ));
   AOI21X1TS U2626 (.Y(n6742), 
	.B0(FE_OFN821_n7619), 
	.A1(n4761), 
	.A0(\fifo_from_fir/fifo_cell1/controller/valid_read ));
   OAI21XLTS U2627 (.Y(n6743), 
	.B0(n4761), 
	.A1(n4763), 
	.A0(\fifo_from_fir/fifo_cell1/data_out/N35 ));
   AOI21X1TS U1995 (.Y(n6213), 
	.B0(FE_OFN791_n7619), 
	.A1(n4575), 
	.A0(\fifo_from_fft/fifo_cell1/controller/valid_read ));
   AO22XLTS U1987 (.Y(n6206), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[6] ), 
	.B0(FE_OFN9_n4574), 
	.A1(FE_OFN1589_acc_fft_data_in_6_), 
	.A0(FE_OFN330_n4573));
   NAND3XLTS U2051 (.Y(n4459), 
	.C(n4640), 
	.B(n4460), 
	.A(FE_OFN327_n4573));
   NAND3XLTS U2682 (.Y(n4645), 
	.C(n4826), 
	.B(n4646), 
	.A(FE_OFN666_n4759));
   OAI21X1TS U3543 (.Y(n3958), 
	.B0(FE_OFN700_n3959), 
	.A1(n5255), 
	.A0(\fifo_to_fft/fifo_cell15/reg_gtok/token ));
   INVXLTS U805 (.Y(n3842), 
	.A(n3844));
   AOI22X1TS U258 (.Y(n3500), 
	.B1(\router/addr_calc/iir_write_calc/counter/N64 ), 
	.B0(FE_OFN932_n3487), 
	.A1(FE_OFN950_n3486), 
	.A0(n7144));
   OAI21XLTS U2701 (.Y(n6761), 
	.B0(n3756), 
	.A1(n7603), 
	.A0(n4830));
   AO22XLTS U2623 (.Y(n6740), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[1] ), 
	.B0(FE_OFN340_n4760), 
	.A1(FE_OFN1804_acc_fir_data_in_1_), 
	.A0(FE_OFN671_n4759));
   AO22XLTS U2624 (.Y(n6741), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[0] ), 
	.B0(FE_OFN338_n4760), 
	.A1(FE_OFN1814_acc_fir_data_in_0_), 
	.A0(FE_OFN671_n4759));
   AO22XLTS U2622 (.Y(n6739), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[2] ), 
	.B0(FE_OFN338_n4760), 
	.A1(FE_OFN1797_acc_fir_data_in_2_), 
	.A0(FE_OFN670_n4759));
   INVX1TS U3523 (.Y(n4001), 
	.A(n3855));
   AO22XLTS U2621 (.Y(n6738), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[3] ), 
	.B0(FE_OFN340_n4760), 
	.A1(FE_OFN1794_acc_fir_data_in_3_), 
	.A0(FE_OFN671_n4759));
   AO22XLTS U2620 (.Y(n6737), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[4] ), 
	.B0(FE_OFN342_n4760), 
	.A1(FE_OFN1789_acc_fir_data_in_4_), 
	.A0(FE_OFN670_n4759));
   AO22XLTS U2619 (.Y(n6736), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[5] ), 
	.B0(FE_OFN342_n4760), 
	.A1(FE_OFN1777_acc_fir_data_in_5_), 
	.A0(FE_OFN668_n4759));
   AO22XLTS U2617 (.Y(n6734), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[7] ), 
	.B0(FE_OFN342_n4760), 
	.A1(FE_OFN1767_acc_fir_data_in_7_), 
	.A0(FE_OFN670_n4759));
   AO22XLTS U2595 (.Y(n6712), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[29] ), 
	.B0(FE_OFN348_n4760), 
	.A1(FE_OFN1645_acc_fir_data_in_29_), 
	.A0(FE_OFN669_n4759));
   AO22XLTS U2594 (.Y(n6711), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[30] ), 
	.B0(FE_OFN348_n4760), 
	.A1(FE_OFN1637_acc_fir_data_in_30_), 
	.A0(FE_OFN669_n4759));
   AO22XLTS U2593 (.Y(n6710), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[31] ), 
	.B0(FE_OFN348_n4760), 
	.A1(FE_OFN1632_acc_fir_data_in_31_), 
	.A0(FE_OFN669_n4759));
   OAI2BB1XLTS U891 (.Y(n5514), 
	.B0(n3958), 
	.A1N(n7973), 
	.A0N(\fifo_to_fft/fifo_cell0/reg_gtok/token ));
   OAI211XLTS U2683 (.Y(n4825), 
	.C0(n9465), 
	.B0(\fifo_from_fir/hang[0] ), 
	.A1(n4827), 
	.A0(n8877));
   AO22XLTS U1989 (.Y(n6208), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[4] ), 
	.B0(FE_OFN9_n4574), 
	.A1(FE_OFN1597_acc_fft_data_in_4_), 
	.A0(FE_OFN330_n4573));
   AO22XLTS U1988 (.Y(n6207), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[5] ), 
	.B0(FE_OFN1_n4574), 
	.A1(FE_OFN1594_acc_fft_data_in_5_), 
	.A0(FE_OFN335_n4573));
   OAI211XLTS U2052 (.Y(n4639), 
	.C0(n9469), 
	.B0(\fifo_from_fft/hang[0] ), 
	.A1(n4641), 
	.A0(n8844));
   AO22XLTS U1991 (.Y(n6210), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[2] ), 
	.B0(FE_OFN0_n4574), 
	.A1(FE_OFN1609_acc_fft_data_in_2_), 
	.A0(FE_OFN336_n4573));
   AO22XLTS U1992 (.Y(n6211), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[1] ), 
	.B0(FE_OFN0_n4574), 
	.A1(FE_OFN1616_acc_fft_data_in_1_), 
	.A0(FE_OFN336_n4573));
   AO22XLTS U1993 (.Y(n6212), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[0] ), 
	.B0(FE_OFN2_n4574), 
	.A1(FE_OFN1622_acc_fft_data_in_0_), 
	.A0(FE_OFN334_n4573));
   AO22XLTS U1986 (.Y(n6205), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[7] ), 
	.B0(FE_OFN0_n4574), 
	.A1(FE_OFN1584_acc_fft_data_in_7_), 
	.A0(FE_OFN337_n4573));
   NAND3XLTS U922 (.Y(n3854), 
	.C(n4000), 
	.B(n3855), 
	.A(n3952));
   NAND3XLTS U1066 (.Y(n4029), 
	.C(n4175), 
	.B(n4030), 
	.A(n4127));
   AO22XLTS U1964 (.Y(n6183), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[29] ), 
	.B0(FE_OFN2_n4574), 
	.A1(FE_OFN1465_acc_fft_data_in_29_), 
	.A0(FE_OFN334_n4573));
   AO22XLTS U1963 (.Y(n6182), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[30] ), 
	.B0(FE_OFN3_n4574), 
	.A1(FE_OFN1458_acc_fft_data_in_30_), 
	.A0(FE_OFN334_n4573));
   AO22XLTS U1962 (.Y(n6181), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[31] ), 
	.B0(FE_OFN3_n4574), 
	.A1(FE_OFN1452_acc_fft_data_in_31_), 
	.A0(FE_OFN333_n4573));
   AO22XLTS U1990 (.Y(n6209), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[3] ), 
	.B0(FE_OFN2_n4574), 
	.A1(FE_OFN1603_acc_fft_data_in_3_), 
	.A0(FE_OFN335_n4573));
   OAI2BB1XLTS U1035 (.Y(n5566), 
	.B0(n4133), 
	.A1N(n7616), 
	.A0N(\fifo_to_fir/fifo_cell0/reg_gtok/token ));
   AOI22X1TS U256 (.Y(n3499), 
	.B1(\router/addr_calc/iir_write_calc/counter/N65 ), 
	.B0(FE_OFN932_n3487), 
	.A1(FE_OFN950_n3486), 
	.A0(FE_OFN1440_router_addr_calc_iir_write_calc_count_19_));
   AO22XLTS U1965 (.Y(n6184), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[28] ), 
	.B0(FE_OFN3_n4574), 
	.A1(FE_OFN1821_acc_fft_data_in_28_), 
	.A0(FE_OFN333_n4573));
   OAI211XLTS U923 (.Y(n3999), 
	.C0(n9477), 
	.B0(\fifo_to_fft/hang[1] ), 
	.A1(n4001), 
	.A0(n8812));
   AO22XLTS U2596 (.Y(n6713), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[28] ), 
	.B0(FE_OFN348_n4760), 
	.A1(FE_OFN1650_acc_fir_data_in_28_), 
	.A0(FE_OFN669_n4759));
   AOI22X1TS U254 (.Y(n3498), 
	.B1(\router/addr_calc/iir_write_calc/counter/N66 ), 
	.B0(FE_OFN931_n3487), 
	.A1(FE_OFN946_n3486), 
	.A0(n7150));
   AO22XLTS U2602 (.Y(n6719), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[22] ), 
	.B0(FE_OFN344_n4760), 
	.A1(FE_OFN1679_acc_fir_data_in_22_), 
	.A0(FE_OFN675_n4759));
   AO22XLTS U2599 (.Y(n6716), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[25] ), 
	.B0(FE_OFN347_n4760), 
	.A1(FE_OFN1665_acc_fir_data_in_25_), 
	.A0(n4759));
   AO22XLTS U2601 (.Y(n6718), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[23] ), 
	.B0(FE_OFN339_n4760), 
	.A1(FE_OFN1675_acc_fir_data_in_23_), 
	.A0(FE_OFN674_n4759));
   AO22XLTS U2603 (.Y(n6720), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[21] ), 
	.B0(FE_OFN344_n4760), 
	.A1(FE_OFN1684_acc_fir_data_in_21_), 
	.A0(FE_OFN675_n4759));
   AO22XLTS U2600 (.Y(n6717), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[24] ), 
	.B0(FE_OFN347_n4760), 
	.A1(FE_OFN1670_acc_fir_data_in_24_), 
	.A0(n4759));
   AO22XLTS U2604 (.Y(n6721), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[20] ), 
	.B0(n4760), 
	.A1(FE_OFN1691_acc_fir_data_in_20_), 
	.A0(FE_OFN672_n4759));
   AO22XLTS U2605 (.Y(n6722), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[19] ), 
	.B0(FE_OFN341_n4760), 
	.A1(FE_OFN1698_acc_fir_data_in_19_), 
	.A0(FE_OFN673_n4759));
   AO22XLTS U2597 (.Y(n6714), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[27] ), 
	.B0(FE_OFN345_n4760), 
	.A1(FE_OFN1655_acc_fir_data_in_27_), 
	.A0(FE_OFN667_n4759));
   AO22XLTS U2606 (.Y(n6723), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[18] ), 
	.B0(FE_OFN346_n4760), 
	.A1(FE_OFN1704_acc_fir_data_in_18_), 
	.A0(FE_OFN676_n4759));
   AO22XLTS U2607 (.Y(n6724), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[17] ), 
	.B0(FE_OFN341_n4760), 
	.A1(FE_OFN1708_acc_fir_data_in_17_), 
	.A0(FE_OFN673_n4759));
   AO22XLTS U2598 (.Y(n6715), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[26] ), 
	.B0(FE_OFN347_n4760), 
	.A1(FE_OFN1658_acc_fir_data_in_26_), 
	.A0(FE_OFN667_n4759));
   AO22XLTS U2609 (.Y(n6726), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[15] ), 
	.B0(FE_OFN339_n4760), 
	.A1(FE_OFN1722_acc_fir_data_in_15_), 
	.A0(FE_OFN674_n4759));
   AO22XLTS U2608 (.Y(n6725), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[16] ), 
	.B0(FE_OFN341_n4760), 
	.A1(FE_OFN1715_acc_fir_data_in_16_), 
	.A0(FE_OFN673_n4759));
   AO22XLTS U2612 (.Y(n6729), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[12] ), 
	.B0(FE_OFN344_n4760), 
	.A1(FE_OFN1737_acc_fir_data_in_12_), 
	.A0(FE_OFN675_n4759));
   AO22XLTS U2613 (.Y(n6730), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[11] ), 
	.B0(FE_OFN346_n4760), 
	.A1(FE_OFN1742_acc_fir_data_in_11_), 
	.A0(FE_OFN677_n4759));
   AO22XLTS U2614 (.Y(n6731), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[10] ), 
	.B0(FE_OFN343_n4760), 
	.A1(FE_OFN1750_acc_fir_data_in_10_), 
	.A0(FE_OFN676_n4759));
   AO22XLTS U2615 (.Y(n6732), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[9] ), 
	.B0(FE_OFN346_n4760), 
	.A1(FE_OFN1753_acc_fir_data_in_9_), 
	.A0(FE_OFN677_n4759));
   AO22XLTS U2616 (.Y(n6733), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[8] ), 
	.B0(FE_OFN346_n4760), 
	.A1(FE_OFN1758_acc_fir_data_in_8_), 
	.A0(FE_OFN677_n4759));
   AO22XLTS U1980 (.Y(n6199), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[13] ), 
	.B0(FE_OFN6_n4574), 
	.A1(FE_OFN1551_acc_fft_data_in_13_), 
	.A0(FE_OFN329_n4573));
   AO22XLTS U1979 (.Y(n6198), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[14] ), 
	.B0(FE_OFN8_n4574), 
	.A1(FE_OFN1546_acc_fft_data_in_14_), 
	.A0(FE_OFN328_n4573));
   AO22XLTS U1978 (.Y(n6197), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[15] ), 
	.B0(FE_OFN7_n4574), 
	.A1(FE_OFN1542_acc_fft_data_in_15_), 
	.A0(FE_OFN329_n4573));
   AO22XLTS U2611 (.Y(n6728), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[13] ), 
	.B0(FE_OFN343_n4760), 
	.A1(FE_OFN1734_acc_fir_data_in_13_), 
	.A0(FE_OFN676_n4759));
   AO22XLTS U2610 (.Y(n6727), 
	.B1(\fifo_from_fir/fifo_cell1/sr_out[14] ), 
	.B0(FE_OFN344_n4760), 
	.A1(FE_OFN1728_acc_fir_data_in_14_), 
	.A0(FE_OFN675_n4759));
   AO22XLTS U1966 (.Y(n6185), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[27] ), 
	.B0(FE_OFN1_n4574), 
	.A1(FE_OFN1473_acc_fft_data_in_27_), 
	.A0(FE_OFN336_n4573));
   AO22XLTS U1977 (.Y(n6196), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[16] ), 
	.B0(FE_OFN9_n4574), 
	.A1(FE_OFN1537_acc_fft_data_in_16_), 
	.A0(FE_OFN327_n4573));
   AO22XLTS U1970 (.Y(n6189), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[23] ), 
	.B0(FE_OFN7_n4574), 
	.A1(FE_OFN1494_acc_fft_data_in_23_), 
	.A0(FE_OFN330_n4573));
   AO22XLTS U1968 (.Y(n6187), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[25] ), 
	.B0(n4574), 
	.A1(FE_OFN1483_acc_fft_data_in_25_), 
	.A0(FE_OFN337_n4573));
   AO22XLTS U1972 (.Y(n6191), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[21] ), 
	.B0(FE_OFN4_n4574), 
	.A1(FE_OFN1505_acc_fft_data_in_21_), 
	.A0(FE_OFN333_n4573));
   AO22XLTS U1971 (.Y(n6190), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[22] ), 
	.B0(FE_OFN4_n4574), 
	.A1(FE_OFN1498_acc_fft_data_in_22_), 
	.A0(FE_OFN332_n4573));
   AO22XLTS U1982 (.Y(n6201), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[11] ), 
	.B0(FE_OFN5_n4574), 
	.A1(FE_OFN1560_acc_fft_data_in_11_), 
	.A0(FE_OFN331_n4573));
   AO22XLTS U1983 (.Y(n6202), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[10] ), 
	.B0(FE_OFN4_n4574), 
	.A1(FE_OFN1564_acc_fft_data_in_10_), 
	.A0(FE_OFN332_n4573));
   AO22XLTS U1985 (.Y(n6204), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[8] ), 
	.B0(FE_OFN5_n4574), 
	.A1(FE_OFN1577_acc_fft_data_in_8_), 
	.A0(FE_OFN332_n4573));
   AO22XLTS U1981 (.Y(n6200), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[12] ), 
	.B0(FE_OFN8_n4574), 
	.A1(FE_OFN1556_acc_fft_data_in_12_), 
	.A0(FE_OFN328_n4573));
   AO22XLTS U1974 (.Y(n6193), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[19] ), 
	.B0(FE_OFN9_n4574), 
	.A1(FE_OFN1515_acc_fft_data_in_19_), 
	.A0(FE_OFN327_n4573));
   AO22XLTS U1973 (.Y(n6192), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[20] ), 
	.B0(FE_OFN6_n4574), 
	.A1(FE_OFN1514_acc_fft_data_in_20_), 
	.A0(FE_OFN331_n4573));
   AO22XLTS U1967 (.Y(n6186), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[26] ), 
	.B0(FE_OFN1_n4574), 
	.A1(FE_OFN1478_acc_fft_data_in_26_), 
	.A0(FE_OFN335_n4573));
   AO22XLTS U1984 (.Y(n6203), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[9] ), 
	.B0(FE_OFN5_n4574), 
	.A1(FE_OFN1572_acc_fft_data_in_9_), 
	.A0(FE_OFN331_n4573));
   AO22XLTS U1976 (.Y(n6195), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[17] ), 
	.B0(FE_OFN8_n4574), 
	.A1(FE_OFN1530_acc_fft_data_in_17_), 
	.A0(FE_OFN328_n4573));
   AO22XLTS U1975 (.Y(n6194), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[18] ), 
	.B0(FE_OFN7_n4574), 
	.A1(FE_OFN1522_acc_fft_data_in_18_), 
	.A0(FE_OFN330_n4573));
   AO22XLTS U1969 (.Y(n6188), 
	.B1(\fifo_from_fft/fifo_cell1/sr_out[24] ), 
	.B0(n4574), 
	.A1(FE_OFN1488_acc_fft_data_in_24_), 
	.A0(FE_OFN337_n4573));
   OAI21XLTS U880 (.Y(n3945), 
	.B0(n3947), 
	.A1(n3943), 
	.A0(n7326));
   AOI22X1TS U477 (.Y(n3629), 
	.B1(\router/addr_calc/fft_write_calc/counter/N67 ), 
	.B0(FE_OFN953_n3619), 
	.A1(FE_OFN971_n3618), 
	.A0(FE_OFN1252_n7397));
   NAND2XLTS U553 (.Y(\router/addr_calc/fft_read_calc/counter/N198 ), 
	.B(n3674), 
	.A(n9439));
   AOI22X1TS U552 (.Y(n3673), 
	.B1(\router/addr_calc/fft_read_calc/counter/N67 ), 
	.B0(FE_OFN874_n3663), 
	.A1(FE_OFN884_n3662), 
	.A0(n7521));
   AOI22X1TS U252 (.Y(n3497), 
	.B1(\router/addr_calc/iir_write_calc/counter/N67 ), 
	.B0(FE_OFN931_n3487), 
	.A1(FE_OFN946_n3486), 
	.A0(n7156));
   AOI21X1TS U1023 (.Y(n5559), 
	.B0(FE_OFN790_n7619), 
	.A1(n4120), 
	.A0(\fifo_to_fir/fifo_cell3/controller/valid_read ));
   OAI21XLTS U1960 (.Y(n4569), 
	.B0(n8472), 
	.A1(n4572), 
	.A0(n7519));
   AOI21X1TS U879 (.Y(n5507), 
	.B0(FE_OFN805_n7619), 
	.A1(n3945), 
	.A0(\fifo_to_fft/fifo_cell3/controller/valid_read ));
   OAI21XLTS U2591 (.Y(n4755), 
	.B0(n8137), 
	.A1(n4758), 
	.A0(n7594));
   NAND3XLTS U1064 (.Y(n4031), 
	.C(n4172), 
	.B(n4032), 
	.A(n4122));
   NAND3XLTS U920 (.Y(n3856), 
	.C(n3997), 
	.B(n3857), 
	.A(n3947));
   OAI21XLTS U877 (.Y(n5506), 
	.B0(n3945), 
	.A1(n3944), 
	.A0(\fifo_to_fft/fifo_cell3/data_out/N35 ));
   AOI22X1TS U562 (.Y(n3678), 
	.B1(\router/addr_calc/fft_read_calc/counter/N62 ), 
	.B0(FE_OFN876_n3663), 
	.A1(FE_OFN886_n3662), 
	.A0(\router/addr_calc/fft_read_calc/count[16] ));
   AOI22X1TS U560 (.Y(n3677), 
	.B1(\router/addr_calc/fft_read_calc/counter/N63 ), 
	.B0(FE_OFN876_n3663), 
	.A1(FE_OFN886_n3662), 
	.A0(n7536));
   AOI22X1TS U558 (.Y(n3676), 
	.B1(\router/addr_calc/fft_read_calc/counter/N64 ), 
	.B0(FE_OFN876_n3663), 
	.A1(FE_OFN884_n3662), 
	.A0(n7531));
   AOI22X1TS U556 (.Y(n3675), 
	.B1(\router/addr_calc/fft_read_calc/counter/N65 ), 
	.B0(FE_OFN876_n3663), 
	.A1(FE_OFN886_n3662), 
	.A0(FE_OFN1258_router_addr_calc_fft_read_calc_count_19_));
   AOI22X1TS U487 (.Y(n3634), 
	.B1(\router/addr_calc/fft_write_calc/counter/N62 ), 
	.B0(FE_OFN956_n3619), 
	.A1(FE_OFN967_n3618), 
	.A0(n7417));
   AOI22X1TS U485 (.Y(n3633), 
	.B1(\router/addr_calc/fft_write_calc/counter/N63 ), 
	.B0(FE_OFN955_n3619), 
	.A1(FE_OFN967_n3618), 
	.A0(n7412));
   AOI22X1TS U483 (.Y(n3632), 
	.B1(\router/addr_calc/fft_write_calc/counter/N64 ), 
	.B0(FE_OFN955_n3619), 
	.A1(FE_OFN968_n3618), 
	.A0(n7407));
   AOI22X1TS U481 (.Y(n3631), 
	.B1(\router/addr_calc/fft_write_calc/counter/N65 ), 
	.B0(FE_OFN953_n3619), 
	.A1(FE_OFN968_n3618), 
	.A0(\router/addr_calc/fft_write_calc/count[19] ));
   AOI22X1TS U250 (.Y(n3496), 
	.B1(\router/addr_calc/iir_write_calc/counter/N68 ), 
	.B0(FE_OFN931_n3487), 
	.A1(FE_OFN946_n3486), 
	.A0(n7162));
   OAI211XLTS U1065 (.Y(n4171), 
	.C0(n9473), 
	.B0(\fifo_to_fir/hang[2] ), 
	.A1(n4173), 
	.A0(n8790));
   OAI211XLTS U921 (.Y(n3996), 
	.C0(n9477), 
	.B0(\fifo_to_fft/hang[2] ), 
	.A1(n3998), 
	.A0(n8811));
   AO22XLTS U2567 (.Y(n6687), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[20] ), 
	.B0(FE_OFN355_n4754), 
	.A1(FE_OFN1694_acc_fir_data_in_20_), 
	.A0(n8143));
   NAND3XLTS U2680 (.Y(n4647), 
	.C(n4823), 
	.B(n4648), 
	.A(n8137));
   NAND3XLTS U2049 (.Y(n4461), 
	.C(n4637), 
	.B(n4462), 
	.A(n8472));
   AO22XLTS U1934 (.Y(n6156), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[22] ), 
	.B0(FE_OFN15_n4568), 
	.A1(FE_OFN1504_acc_fft_data_in_22_), 
	.A0(n8478));
   AOI21X1TS U2589 (.Y(n6708), 
	.B0(FE_OFN809_n7619), 
	.A1(n4755), 
	.A0(\fifo_from_fir/fifo_cell2/controller/valid_read ));
   OAI21XLTS U1959 (.Y(n6180), 
	.B0(n4569), 
	.A1(n4571), 
	.A0(\fifo_from_fft/fifo_cell2/data_out/N35 ));
   OAI21XLTS U2590 (.Y(n6709), 
	.B0(n4755), 
	.A1(n4757), 
	.A0(\fifo_from_fir/fifo_cell2/data_out/N35 ));
   AOI21X1TS U1958 (.Y(n6179), 
	.B0(FE_OFN807_n7619), 
	.A1(n4569), 
	.A0(\fifo_from_fft/fifo_cell2/controller/valid_read ));
   AOI22X1TS U495 (.Y(n3638), 
	.B1(\router/addr_calc/fft_write_calc/counter/N58 ), 
	.B0(FE_OFN956_n3619), 
	.A1(FE_OFN967_n3618), 
	.A0(n7432));
   AOI22X1TS U248 (.Y(n3495), 
	.B1(\router/addr_calc/iir_write_calc/counter/N69 ), 
	.B0(n3487), 
	.A1(FE_OFN944_n3486), 
	.A0(FE_OFN1244_router_addr_calc_iir_write_calc_count_23_));
   AOI22X1TS U582 (.Y(n3688), 
	.B1(\router/addr_calc/fft_read_calc/counter/N52 ), 
	.B0(FE_OFN867_n3663), 
	.A1(FE_OFN882_n3662), 
	.A0(n7581));
   AOI22X1TS U580 (.Y(n3687), 
	.B1(\router/addr_calc/fft_read_calc/counter/N53 ), 
	.B0(FE_OFN867_n3663), 
	.A1(FE_OFN882_n3662), 
	.A0(n7576));
   AOI22X1TS U327 (.Y(n3541), 
	.B1(\router/addr_calc/fir_write_calc/counter/N67 ), 
	.B0(FE_OFN891_n3531), 
	.A1(FE_OFN902_n3530), 
	.A0(FE_OFN1254_n7159));
   AOI22X1TS U511 (.Y(n3646), 
	.B1(\router/addr_calc/fft_write_calc/counter/N50 ), 
	.B0(FE_OFN960_n3619), 
	.A1(FE_OFN963_n3618), 
	.A0(n7467));
   AOI22X1TS U568 (.Y(n3681), 
	.B1(\router/addr_calc/fft_read_calc/counter/N59 ), 
	.B0(FE_OFN871_n3663), 
	.A1(FE_OFN887_n3662), 
	.A0(n7551));
   AOI22X1TS U493 (.Y(n3637), 
	.B1(\router/addr_calc/fft_write_calc/counter/N59 ), 
	.B0(FE_OFN957_n3619), 
	.A1(FE_OFN966_n3618), 
	.A0(n7427));
   AOI22X1TS U505 (.Y(n3643), 
	.B1(\router/addr_calc/fft_write_calc/counter/N53 ), 
	.B0(FE_OFN959_n3619), 
	.A1(FE_OFN964_n3618), 
	.A0(n7452));
   NAND2XLTS U549 (.Y(\router/addr_calc/fft_read_calc/counter/N200 ), 
	.B(n3672), 
	.A(n9439));
   AOI22X1TS U503 (.Y(n3642), 
	.B1(\router/addr_calc/fft_write_calc/counter/N54 ), 
	.B0(FE_OFN958_n3619), 
	.A1(FE_OFN964_n3618), 
	.A0(n7447));
   AOI22X1TS U566 (.Y(n3680), 
	.B1(\router/addr_calc/fft_read_calc/counter/N60 ), 
	.B0(FE_OFN871_n3663), 
	.A1(FE_OFN887_n3662), 
	.A0(n7546));
   AOI22X1TS U584 (.Y(n3689), 
	.B1(\router/addr_calc/fft_read_calc/counter/N51 ), 
	.B0(FE_OFN868_n3663), 
	.A1(FE_OFN881_n3662), 
	.A0(\router/addr_calc/fft_read_calc/count[5] ));
   AOI22X1TS U473 (.Y(n3627), 
	.B1(\router/addr_calc/fft_write_calc/counter/N69 ), 
	.B0(FE_OFN951_n3619), 
	.A1(FE_OFN969_n3618), 
	.A0(\router/addr_calc/fft_write_calc/count[23] ));
   AOI22X1TS U586 (.Y(n3690), 
	.B1(\router/addr_calc/fft_read_calc/counter/N50 ), 
	.B0(FE_OFN875_n3663), 
	.A1(FE_OFN877_n3662), 
	.A0(n7586));
   AOI22X1TS U548 (.Y(n3671), 
	.B1(\router/addr_calc/fft_read_calc/counter/N69 ), 
	.B0(FE_OFN872_n3663), 
	.A1(FE_OFN883_n3662), 
	.A0(\router/addr_calc/fft_read_calc/count[23] ));
   AOI22X1TS U398 (.Y(n3583), 
	.B1(\router/addr_calc/fir_read_calc/counter/N69 ), 
	.B0(FE_OFN916_n3575), 
	.A1(FE_OFN927_n3574), 
	.A0(\router/addr_calc/fir_read_calc/count[23] ));
   AOI22X1TS U491 (.Y(n3636), 
	.B1(\router/addr_calc/fft_write_calc/counter/N60 ), 
	.B0(FE_OFN956_n3619), 
	.A1(FE_OFN966_n3618), 
	.A0(n7422));
   AOI22X1TS U513 (.Y(n3647), 
	.B1(\router/addr_calc/fft_write_calc/counter/N49 ), 
	.B0(FE_OFN960_n3619), 
	.A1(FE_OFN963_n3618), 
	.A0(n7472));
   AOI22X1TS U570 (.Y(n3682), 
	.B1(\router/addr_calc/fft_read_calc/counter/N58 ), 
	.B0(FE_OFN871_n3663), 
	.A1(FE_OFN887_n3662), 
	.A0(n7556));
   AOI22X1TS U588 (.Y(n3691), 
	.B1(\router/addr_calc/fft_read_calc/counter/N49 ), 
	.B0(FE_OFN875_n3663), 
	.A1(n3662), 
	.A0(n7591));
   AOI22X1TS U574 (.Y(n3684), 
	.B1(\router/addr_calc/fft_read_calc/counter/N56 ), 
	.B0(FE_OFN869_n3663), 
	.A1(FE_OFN885_n3662), 
	.A0(n7566));
   AOI22X1TS U592 (.Y(n3693), 
	.B1(\router/addr_calc/fft_read_calc/counter/N47 ), 
	.B0(FE_OFN873_n3663), 
	.A1(FE_OFN877_n3662), 
	.A0(n7601));
   AOI22X1TS U402 (.Y(n3585), 
	.B1(\router/addr_calc/fir_read_calc/counter/N67 ), 
	.B0(FE_OFN916_n3575), 
	.A1(FE_OFN926_n3574), 
	.A0(FE_OFN1253_n7283));
   AOI22X1TS U507 (.Y(n3644), 
	.B1(\router/addr_calc/fft_write_calc/counter/N52 ), 
	.B0(FE_OFN959_n3619), 
	.A1(FE_OFN962_n3618), 
	.A0(n7457));
   AOI22X1TS U578 (.Y(n3686), 
	.B1(\router/addr_calc/fft_read_calc/counter/N54 ), 
	.B0(FE_OFN869_n3663), 
	.A1(FE_OFN882_n3662), 
	.A0(n7571));
   AOI22X1TS U499 (.Y(n3640), 
	.B1(\router/addr_calc/fft_write_calc/counter/N56 ), 
	.B0(FE_OFN958_n3619), 
	.A1(FE_OFN965_n3618), 
	.A0(n7442));
   AOI22X1TS U590 (.Y(n3692), 
	.B1(\router/addr_calc/fft_read_calc/counter/N48 ), 
	.B0(FE_OFN875_n3663), 
	.A1(n3662), 
	.A0(n7596));
   AOI22X1TS U515 (.Y(n3648), 
	.B1(\router/addr_calc/fft_write_calc/counter/N48 ), 
	.B0(FE_OFN960_n3619), 
	.A1(FE_OFN963_n3618), 
	.A0(n7477));
   AOI22X1TS U564 (.Y(n3679), 
	.B1(\router/addr_calc/fft_read_calc/counter/N61 ), 
	.B0(FE_OFN871_n3663), 
	.A1(FE_OFN887_n3662), 
	.A0(n7541));
   AOI22X1TS U594 (.Y(n3694), 
	.B1(n7957), 
	.B0(FE_OFN873_n3663), 
	.A1(FE_OFN878_n3662), 
	.A0(\router/addr_calc/fft_read_calc/count[0] ));
   AOI22X1TS U489 (.Y(n3635), 
	.B1(\router/addr_calc/fft_write_calc/counter/N61 ), 
	.B0(FE_OFN957_n3619), 
	.A1(FE_OFN966_n3618), 
	.A0(FE_OFN1270_router_addr_calc_fft_write_calc_count_15_));
   AOI22X1TS U517 (.Y(n3649), 
	.B1(\router/addr_calc/fft_write_calc/counter/N47 ), 
	.B0(n3619), 
	.A1(FE_OFN970_n3618), 
	.A0(n7482));
   AOI22X1TS U519 (.Y(n3650), 
	.B1(n7958), 
	.B0(n3619), 
	.A1(FE_OFN970_n3618), 
	.A0(\router/addr_calc/fft_write_calc/count[0] ));
   AOI22X1TS U509 (.Y(n3645), 
	.B1(\router/addr_calc/fft_write_calc/counter/N51 ), 
	.B0(FE_OFN959_n3619), 
	.A1(FE_OFN962_n3618), 
	.A0(n7462));
   AOI22X1TS U323 (.Y(n3539), 
	.B1(\router/addr_calc/fir_write_calc/counter/N69 ), 
	.B0(FE_OFN891_n3531), 
	.A1(FE_OFN902_n3530), 
	.A0(FE_OFN1248_router_addr_calc_fir_write_calc_count_23_));
   AO22XLTS U1933 (.Y(n6155), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[23] ), 
	.B0(FE_OFN15_n4568), 
	.A1(FE_OFN1495_acc_fft_data_in_23_), 
	.A0(n8478));
   OAI21XLTS U1019 (.Y(n4115), 
	.B0(n4117), 
	.A1(n4113), 
	.A0(n7430));
   OAI211XLTS U2681 (.Y(n4822), 
	.C0(n9466), 
	.B0(\fifo_from_fir/hang[1] ), 
	.A1(n4824), 
	.A0(n8877));
   AO22XLTS U1935 (.Y(n6157), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[21] ), 
	.B0(FE_OFN16_n4568), 
	.A1(FE_OFN1508_acc_fft_data_in_21_), 
	.A0(n8478));
   AO22XLTS U1926 (.Y(n6148), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[30] ), 
	.B0(FE_OFN18_n4568), 
	.A1(FE_OFN1462_acc_fft_data_in_30_), 
	.A0(n8480));
   AO22XLTS U1936 (.Y(n6158), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[20] ), 
	.B0(FE_OFN15_n4568), 
	.A1(FE_OFN1513_acc_fft_data_in_20_), 
	.A0(n8478));
   AO22XLTS U1940 (.Y(n6162), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[16] ), 
	.B0(n4568), 
	.A1(FE_OFN1534_acc_fft_data_in_16_), 
	.A0(n8477));
   AO22XLTS U1937 (.Y(n6159), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[19] ), 
	.B0(FE_OFN10_n4568), 
	.A1(FE_OFN1515_acc_fft_data_in_19_), 
	.A0(n8477));
   AO22XLTS U1939 (.Y(n6161), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[17] ), 
	.B0(n4568), 
	.A1(FE_OFN1532_acc_fft_data_in_17_), 
	.A0(n8477));
   AO22XLTS U1938 (.Y(n6160), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[18] ), 
	.B0(FE_OFN10_n4568), 
	.A1(FE_OFN1526_acc_fft_data_in_18_), 
	.A0(n8477));
   AO22XLTS U1925 (.Y(n6147), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[31] ), 
	.B0(FE_OFN16_n4568), 
	.A1(FE_OFN1456_acc_fft_data_in_31_), 
	.A0(n8480));
   AO22XLTS U2565 (.Y(n6685), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[22] ), 
	.B0(FE_OFN356_n4754), 
	.A1(FE_OFN1679_acc_fir_data_in_22_), 
	.A0(n8143));
   AO22XLTS U1927 (.Y(n6149), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[29] ), 
	.B0(FE_OFN17_n4568), 
	.A1(FE_OFN1467_acc_fft_data_in_29_), 
	.A0(n8480));
   OAI21XLTS U875 (.Y(n3940), 
	.B0(n3942), 
	.A1(n3938), 
	.A0(n7321));
   AO22XLTS U2564 (.Y(n6684), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[23] ), 
	.B0(FE_OFN355_n4754), 
	.A1(FE_OFN1677_acc_fir_data_in_23_), 
	.A0(n8143));
   AO22XLTS U2566 (.Y(n6686), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[21] ), 
	.B0(FE_OFN356_n4754), 
	.A1(FE_OFN1685_acc_fir_data_in_21_), 
	.A0(n8143));
   AO22XLTS U2559 (.Y(n6679), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[28] ), 
	.B0(FE_OFN353_n4754), 
	.A1(FE_OFN1648_acc_fir_data_in_28_), 
	.A0(n8145));
   OAI211XLTS U2050 (.Y(n4636), 
	.C0(n9469), 
	.B0(\fifo_from_fft/hang[1] ), 
	.A1(n4638), 
	.A0(n8844));
   NAND2XLTS U496 (.Y(\router/addr_calc/fft_write_calc/counter/N189 ), 
	.B(n3639), 
	.A(n9445));
   NAND2XLTS U571 (.Y(\router/addr_calc/fft_read_calc/counter/N189 ), 
	.B(n3683), 
	.A(n9436));
   NAND2XLTS U500 (.Y(\router/addr_calc/fft_write_calc/counter/N187 ), 
	.B(n3641), 
	.A(n9444));
   AOI22X1TS U408 (.Y(n3588), 
	.B1(\router/addr_calc/fir_read_calc/counter/N64 ), 
	.B0(FE_OFN915_n3575), 
	.A1(FE_OFN925_n3574), 
	.A0(n7293));
   AOI22X1TS U406 (.Y(n3587), 
	.B1(\router/addr_calc/fir_read_calc/counter/N65 ), 
	.B0(FE_OFN915_n3575), 
	.A1(FE_OFN926_n3574), 
	.A0(\router/addr_calc/fir_read_calc/count[19] ));
   AOI22X1TS U410 (.Y(n3589), 
	.B1(\router/addr_calc/fir_read_calc/counter/N63 ), 
	.B0(FE_OFN914_n3575), 
	.A1(FE_OFN925_n3574), 
	.A0(FE_OFN1262_n7298));
   AOI22X1TS U337 (.Y(n3546), 
	.B1(\router/addr_calc/fir_write_calc/counter/N62 ), 
	.B0(FE_OFN896_n3531), 
	.A1(FE_OFN908_n3530), 
	.A0(\router/addr_calc/fir_write_calc/count[16] ));
   AOI22X1TS U396 (.Y(n3582), 
	.B1(\router/addr_calc/fir_read_calc/counter/N70 ), 
	.B0(FE_OFN917_n3575), 
	.A1(FE_OFN927_n3574), 
	.A0(FE_OFN1243_n7273));
   AOI22X1TS U246 (.Y(n3494), 
	.B1(\router/addr_calc/iir_write_calc/counter/N70 ), 
	.B0(FE_OFN930_n3487), 
	.A1(FE_OFN944_n3486), 
	.A0(n7168));
   AOI22X1TS U333 (.Y(n3544), 
	.B1(\router/addr_calc/fir_write_calc/counter/N64 ), 
	.B0(FE_OFN895_n3531), 
	.A1(FE_OFN908_n3530), 
	.A0(n7171));
   AOI22X1TS U546 (.Y(n3670), 
	.B1(\router/addr_calc/fft_read_calc/counter/N70 ), 
	.B0(FE_OFN872_n3663), 
	.A1(FE_OFN883_n3662), 
	.A0(n7511));
   AOI22X1TS U471 (.Y(n3626), 
	.B1(\router/addr_calc/fft_write_calc/counter/N70 ), 
	.B0(FE_OFN951_n3619), 
	.A1(FE_OFN970_n3618), 
	.A0(n7387));
   AOI22X1TS U321 (.Y(n3538), 
	.B1(\router/addr_calc/fir_write_calc/counter/N70 ), 
	.B0(FE_OFN893_n3531), 
	.A1(FE_OFN902_n3530), 
	.A0(n7147));
   NAND2XLTS U575 (.Y(\router/addr_calc/fft_read_calc/counter/N187 ), 
	.B(n3685), 
	.A(n9436));
   AOI22X1TS U412 (.Y(n3590), 
	.B1(\router/addr_calc/fir_read_calc/counter/N62 ), 
	.B0(FE_OFN913_n3575), 
	.A1(FE_OFN924_n3574), 
	.A0(FE_OFN1265_n7303));
   AOI22X1TS U335 (.Y(n3545), 
	.B1(\router/addr_calc/fir_write_calc/counter/N63 ), 
	.B0(FE_OFN896_n3531), 
	.A1(FE_OFN908_n3530), 
	.A0(n7177));
   AOI22X1TS U331 (.Y(n3543), 
	.B1(\router/addr_calc/fir_write_calc/counter/N65 ), 
	.B0(FE_OFN895_n3531), 
	.A1(FE_OFN905_n3530), 
	.A0(FE_OFN1261_router_addr_calc_fir_write_calc_count_19_));
   AO22XLTS U2569 (.Y(n6689), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[18] ), 
	.B0(FE_OFN355_n4754), 
	.A1(FE_OFN1706_acc_fir_data_in_18_), 
	.A0(n8142));
   AO22XLTS U2568 (.Y(n6688), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[19] ), 
	.B0(FE_OFN354_n4754), 
	.A1(FE_OFN1697_acc_fir_data_in_19_), 
	.A0(n8142));
   AO22XLTS U2570 (.Y(n6690), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[17] ), 
	.B0(FE_OFN354_n4754), 
	.A1(FE_OFN1711_acc_fir_data_in_17_), 
	.A0(n8142));
   AO22XLTS U2571 (.Y(n6691), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[16] ), 
	.B0(FE_OFN354_n4754), 
	.A1(FE_OFN1718_acc_fir_data_in_16_), 
	.A0(n8142));
   OAI21XLTS U1016 (.Y(n5555), 
	.B0(n4115), 
	.A1(n4114), 
	.A0(\fifo_to_fir/fifo_cell4/data_out/N35 ));
   AO22XLTS U2572 (.Y(n6692), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[15] ), 
	.B0(FE_OFN357_n4754), 
	.A1(FE_OFN1721_acc_fir_data_in_15_), 
	.A0(n8141));
   AO22XLTS U2573 (.Y(n6693), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[14] ), 
	.B0(FE_OFN357_n4754), 
	.A1(FE_OFN1729_acc_fir_data_in_14_), 
	.A0(n8141));
   AO22XLTS U2574 (.Y(n6694), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[13] ), 
	.B0(FE_OFN357_n4754), 
	.A1(FE_OFN1735_acc_fir_data_in_13_), 
	.A0(n8141));
   AO22XLTS U2575 (.Y(n6695), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[12] ), 
	.B0(FE_OFN356_n4754), 
	.A1(FE_OFN1740_acc_fir_data_in_12_), 
	.A0(n8141));
   AO22XLTS U2576 (.Y(n6696), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[11] ), 
	.B0(FE_OFN358_n4754), 
	.A1(FE_OFN1743_acc_fir_data_in_11_), 
	.A0(n8140));
   AO22XLTS U2577 (.Y(n6697), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[10] ), 
	.B0(FE_OFN358_n4754), 
	.A1(FE_OFN1748_acc_fir_data_in_10_), 
	.A0(n8140));
   AO22XLTS U2578 (.Y(n6698), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[9] ), 
	.B0(FE_OFN358_n4754), 
	.A1(FE_OFN1755_acc_fir_data_in_9_), 
	.A0(n8140));
   AO22XLTS U2579 (.Y(n6699), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[8] ), 
	.B0(FE_OFN358_n4754), 
	.A1(FE_OFN1760_acc_fir_data_in_8_), 
	.A0(n8140));
   AO22XLTS U2580 (.Y(n6700), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[7] ), 
	.B0(FE_OFN349_n4754), 
	.A1(FE_OFN1767_acc_fir_data_in_7_), 
	.A0(n8139));
   AO22XLTS U2581 (.Y(n6701), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[6] ), 
	.B0(FE_OFN349_n4754), 
	.A1(FE_OFN1776_acc_fir_data_in_6_), 
	.A0(n8139));
   AO22XLTS U2582 (.Y(n6702), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[5] ), 
	.B0(FE_OFN351_n4754), 
	.A1(FE_OFN1779_acc_fir_data_in_5_), 
	.A0(n8139));
   AO22XLTS U2583 (.Y(n6703), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[4] ), 
	.B0(FE_OFN351_n4754), 
	.A1(FE_OFN1789_acc_fir_data_in_4_), 
	.A0(n8139));
   AO22XLTS U2584 (.Y(n6704), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[3] ), 
	.B0(FE_OFN352_n4754), 
	.A1(FE_OFN1792_acc_fir_data_in_3_), 
	.A0(n8138));
   AO22XLTS U2585 (.Y(n6705), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[2] ), 
	.B0(FE_OFN352_n4754), 
	.A1(FE_OFN1799_acc_fir_data_in_2_), 
	.A0(n8138));
   AO22XLTS U2586 (.Y(n6706), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[1] ), 
	.B0(FE_OFN351_n4754), 
	.A1(FE_OFN1804_acc_fir_data_in_1_), 
	.A0(n8138));
   AO22XLTS U2587 (.Y(n6707), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[0] ), 
	.B0(FE_OFN352_n4754), 
	.A1(FE_OFN1814_acc_fir_data_in_0_), 
	.A0(n8138));
   NAND3XLTS U1062 (.Y(n4033), 
	.C(n4169), 
	.B(n4034), 
	.A(n4117));
   AOI21X1TS U1018 (.Y(n5556), 
	.B0(FE_OFN804_n7619), 
	.A1(n4115), 
	.A0(\fifo_to_fir/fifo_cell4/controller/valid_read ));
   AO22XLTS U1928 (.Y(n6150), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[28] ), 
	.B0(FE_OFN17_n4568), 
	.A1(FE_OFN1471_acc_fft_data_in_28_), 
	.A0(n8480));
   AOI21X1TS U874 (.Y(n5504), 
	.B0(FE_OFN819_n7619), 
	.A1(n3940), 
	.A0(\fifo_to_fft/fifo_cell4/controller/valid_read ));
   OAI21XLTS U872 (.Y(n5503), 
	.B0(n3940), 
	.A1(n3939), 
	.A0(\fifo_to_fft/fifo_cell4/data_out/N35 ));
   NAND3XLTS U918 (.Y(n3858), 
	.C(n3994), 
	.B(n3859), 
	.A(n3942));
   AO22XLTS U2556 (.Y(n6676), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[31] ), 
	.B0(FE_OFN353_n4754), 
	.A1(FE_OFN1631_acc_fir_data_in_31_), 
	.A0(n8145));
   AO22XLTS U2557 (.Y(n6677), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[30] ), 
	.B0(FE_OFN353_n4754), 
	.A1(FE_OFN1634_acc_fir_data_in_30_), 
	.A0(n8145));
   AO22XLTS U2558 (.Y(n6678), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[29] ), 
	.B0(FE_OFN353_n4754), 
	.A1(FE_OFN1644_acc_fir_data_in_29_), 
	.A0(n8145));
   AOI22X1TS U544 (.Y(n3669), 
	.B1(\router/addr_calc/fft_read_calc/counter/N71 ), 
	.B0(n3663), 
	.A1(FE_OFN880_n3662), 
	.A0(n7506));
   AOI22X1TS U394 (.Y(n3581), 
	.B1(\router/addr_calc/fir_read_calc/counter/N71 ), 
	.B0(n3575), 
	.A1(FE_OFN921_n3574), 
	.A0(FE_OFN1242_n7268));
   AOI22X1TS U416 (.Y(n3592), 
	.B1(\router/addr_calc/fir_read_calc/counter/N60 ), 
	.B0(FE_OFN914_n3575), 
	.A1(FE_OFN925_n3574), 
	.A0(FE_OFN1277_n7308));
   AOI22X1TS U343 (.Y(n3549), 
	.B1(\router/addr_calc/fir_write_calc/counter/N59 ), 
	.B0(FE_OFN892_n3531), 
	.A1(FE_OFN907_n3530), 
	.A0(n7195));
   AOI22X1TS U365 (.Y(n3560), 
	.B1(\router/addr_calc/fir_write_calc/counter/N48 ), 
	.B0(FE_OFN888_n3531), 
	.A1(FE_OFN901_n3530), 
	.A0(n7239));
   AOI22X1TS U244 (.Y(n3493), 
	.B1(\router/addr_calc/iir_write_calc/counter/N71 ), 
	.B0(FE_OFN930_n3487), 
	.A1(FE_OFN943_n3486), 
	.A0(n7174));
   AOI22X1TS U424 (.Y(n3596), 
	.B1(\router/addr_calc/fir_read_calc/counter/N56 ), 
	.B0(FE_OFN912_n3575), 
	.A1(FE_OFN923_n3574), 
	.A0(FE_OFN1279_n7328));
   AOI22X1TS U367 (.Y(n3561), 
	.B1(\router/addr_calc/fir_write_calc/counter/N47 ), 
	.B0(n3531), 
	.A1(FE_OFN903_n3530), 
	.A0(n7244));
   AOI22X1TS U341 (.Y(n3548), 
	.B1(\router/addr_calc/fir_write_calc/counter/N60 ), 
	.B0(FE_OFN892_n3531), 
	.A1(FE_OFN907_n3530), 
	.A0(n7189));
   AOI22X1TS U339 (.Y(n3547), 
	.B1(\router/addr_calc/fir_write_calc/counter/N61 ), 
	.B0(FE_OFN896_n3531), 
	.A1(FE_OFN908_n3530), 
	.A0(n7183));
   AOI22X1TS U353 (.Y(n3554), 
	.B1(\router/addr_calc/fir_write_calc/counter/N54 ), 
	.B0(FE_OFN890_n3531), 
	.A1(FE_OFN906_n3530), 
	.A0(n7214));
   CLKINVX1TS U663 (.Y(n5375), 
	.A(n3746));
   AOI22X1TS U430 (.Y(n3599), 
	.B1(\router/addr_calc/fir_read_calc/counter/N53 ), 
	.B0(FE_OFN911_n3575), 
	.A1(FE_OFN922_n3574), 
	.A0(n7338));
   CLKINVX1TS U665 (.Y(n5376), 
	.A(n3747));
   CLKINVX1TS U667 (.Y(n5377), 
	.A(n3748));
   CLKINVX1TS U669 (.Y(n5378), 
	.A(n3749));
   CLKINVX1TS U645 (.Y(n5366), 
	.A(n3737));
   AOI22X1TS U428 (.Y(n3598), 
	.B1(\router/addr_calc/fir_read_calc/counter/N54 ), 
	.B0(FE_OFN911_n3575), 
	.A1(FE_OFN922_n3574), 
	.A0(FE_OFN1278_n7333));
   CLKINVX1TS U671 (.Y(n5379), 
	.A(n3750));
   AOI22X1TS U349 (.Y(n3552), 
	.B1(\router/addr_calc/fir_write_calc/counter/N56 ), 
	.B0(FE_OFN889_n3531), 
	.A1(FE_OFN904_n3530), 
	.A0(n7209));
   CLKINVX1TS U673 (.Y(n5380), 
	.A(n3751));
   CLKINVX1TS U675 (.Y(n5381), 
	.A(n3752));
   AOI22X1TS U432 (.Y(n3600), 
	.B1(\router/addr_calc/fir_read_calc/counter/N52 ), 
	.B0(FE_OFN911_n3575), 
	.A1(FE_OFN920_n3574), 
	.A0(n7343));
   CLKINVX1TS U677 (.Y(n5382), 
	.A(n3753));
   CLKINVX1TS U643 (.Y(n5365), 
	.A(n3736));
   AOI22X1TS U359 (.Y(n3557), 
	.B1(\router/addr_calc/fir_write_calc/counter/N51 ), 
	.B0(FE_OFN897_n3531), 
	.A1(FE_OFN898_n3530), 
	.A0(\router/addr_calc/fir_write_calc/count[5] ));
   CLKINVX1TS U641 (.Y(n5364), 
	.A(n3735));
   AOI22X1TS U369 (.Y(n3562), 
	.B1(n7956), 
	.B0(FE_OFN897_n3531), 
	.A1(FE_OFN898_n3530), 
	.A0(\router/addr_calc/fir_write_calc/count[0] ));
   AOI22X1TS U357 (.Y(n3556), 
	.B1(\router/addr_calc/fir_write_calc/counter/N52 ), 
	.B0(FE_OFN890_n3531), 
	.A1(FE_OFN906_n3530), 
	.A0(n7224));
   AOI22X1TS U469 (.Y(n3625), 
	.B1(\router/addr_calc/fft_write_calc/counter/N71 ), 
	.B0(FE_OFN954_n3619), 
	.A1(FE_OFN971_n3618), 
	.A0(n7382));
   AOI22X1TS U434 (.Y(n3601), 
	.B1(\router/addr_calc/fir_read_calc/counter/N51 ), 
	.B0(FE_OFN910_n3575), 
	.A1(FE_OFN920_n3574), 
	.A0(FE_OFN1276_router_addr_calc_fir_read_calc_count_5_));
   CLKINVX1TS U639 (.Y(n5363), 
	.A(n3734));
   AOI22X1TS U436 (.Y(n3602), 
	.B1(\router/addr_calc/fir_read_calc/counter/N50 ), 
	.B0(FE_OFN909_n3575), 
	.A1(FE_OFN919_n3574), 
	.A0(n7348));
   AOI22X1TS U361 (.Y(n3558), 
	.B1(\router/addr_calc/fir_write_calc/counter/N50 ), 
	.B0(FE_OFN888_n3531), 
	.A1(FE_OFN899_n3530), 
	.A0(n7229));
   AOI22X1TS U420 (.Y(n3594), 
	.B1(\router/addr_calc/fir_read_calc/counter/N58 ), 
	.B0(FE_OFN912_n3575), 
	.A1(FE_OFN923_n3574), 
	.A0(n7318));
   AOI22X1TS U438 (.Y(n3603), 
	.B1(\router/addr_calc/fir_read_calc/counter/N49 ), 
	.B0(FE_OFN909_n3575), 
	.A1(FE_OFN919_n3574), 
	.A0(FE_OFN1275_n7353));
   CLKINVX1TS U637 (.Y(n5362), 
	.A(n3733));
   AOI22X1TS U440 (.Y(n3604), 
	.B1(\router/addr_calc/fir_read_calc/counter/N48 ), 
	.B0(FE_OFN909_n3575), 
	.A1(n3574), 
	.A0(FE_OFN1274_n7358));
   AOI22X1TS U442 (.Y(n3605), 
	.B1(\router/addr_calc/fir_read_calc/counter/N47 ), 
	.B0(n3575), 
	.A1(FE_OFN921_n3574), 
	.A0(n7363));
   CLKINVX1TS U635 (.Y(n5361), 
	.A(n3732));
   AOI22X1TS U444 (.Y(n3606), 
	.B1(n7955), 
	.B0(FE_OFN910_n3575), 
	.A1(FE_OFN922_n3574), 
	.A0(FE_OFN1446_router_addr_calc_fir_read_calc_count_0_));
   AOI22X1TS U414 (.Y(n3591), 
	.B1(\router/addr_calc/fir_read_calc/counter/N61 ), 
	.B0(FE_OFN913_n3575), 
	.A1(FE_OFN924_n3574), 
	.A0(FE_OFN1271_router_addr_calc_fir_read_calc_count_15_));
   CLKINVX1TS U633 (.Y(n5360), 
	.A(n3731));
   AOI22X1TS U319 (.Y(n3537), 
	.B1(\router/addr_calc/fir_write_calc/counter/N71 ), 
	.B0(FE_OFN893_n3531), 
	.A1(FE_OFN900_n3530), 
	.A0(n7141));
   CLKINVX1TS U631 (.Y(n5359), 
	.A(n3730));
   AOI22X1TS U355 (.Y(n3555), 
	.B1(\router/addr_calc/fir_write_calc/counter/N53 ), 
	.B0(FE_OFN890_n3531), 
	.A1(FE_OFN906_n3530), 
	.A0(n7219));
   AOI22X1TS U345 (.Y(n3550), 
	.B1(\router/addr_calc/fir_write_calc/counter/N58 ), 
	.B0(FE_OFN892_n3531), 
	.A1(FE_OFN907_n3530), 
	.A0(n7201));
   AOI22X1TS U363 (.Y(n3559), 
	.B1(\router/addr_calc/fir_write_calc/counter/N49 ), 
	.B0(n3531), 
	.A1(FE_OFN901_n3530), 
	.A0(n7234));
   AOI22X1TS U418 (.Y(n3593), 
	.B1(\router/addr_calc/fir_read_calc/counter/N59 ), 
	.B0(FE_OFN913_n3575), 
	.A1(FE_OFN924_n3574), 
	.A0(n7313));
   AO22XLTS U2562 (.Y(n6682), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[25] ), 
	.B0(n4754), 
	.A1(FE_OFN1661_acc_fir_data_in_25_), 
	.A0(n8144));
   AO22XLTS U2561 (.Y(n6681), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[26] ), 
	.B0(FE_OFN350_n4754), 
	.A1(FE_OFN1659_acc_fir_data_in_26_), 
	.A0(n8144));
   AO22XLTS U2560 (.Y(n6680), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[27] ), 
	.B0(FE_OFN350_n4754), 
	.A1(FE_OFN1654_acc_fir_data_in_27_), 
	.A0(n8144));
   AO22XLTS U2563 (.Y(n6683), 
	.B1(\fifo_from_fir/fifo_cell2/sr_out[24] ), 
	.B0(FE_OFN350_n4754), 
	.A1(FE_OFN1666_acc_fir_data_in_24_), 
	.A0(n8144));
   AO22XLTS U1929 (.Y(n6151), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[27] ), 
	.B0(FE_OFN20_n4568), 
	.A1(FE_OFN1475_acc_fft_data_in_27_), 
	.A0(n8479));
   AO22XLTS U1930 (.Y(n6152), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[26] ), 
	.B0(FE_OFN20_n4568), 
	.A1(FE_OFN1481_acc_fft_data_in_26_), 
	.A0(n8479));
   AO22XLTS U1931 (.Y(n6153), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[25] ), 
	.B0(FE_OFN21_n4568), 
	.A1(FE_OFN1486_acc_fft_data_in_25_), 
	.A0(n8479));
   AO22XLTS U1932 (.Y(n6154), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[24] ), 
	.B0(FE_OFN21_n4568), 
	.A1(FE_OFN1492_acc_fft_data_in_24_), 
	.A0(n8479));
   AO22XLTS U1949 (.Y(n6171), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[7] ), 
	.B0(FE_OFN19_n4568), 
	.A1(FE_OFN1580_acc_fft_data_in_7_), 
	.A0(n8474));
   AO22XLTS U1950 (.Y(n6172), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[6] ), 
	.B0(FE_OFN19_n4568), 
	.A1(FE_OFN1589_acc_fft_data_in_6_), 
	.A0(n8474));
   AO22XLTS U1956 (.Y(n6178), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[0] ), 
	.B0(FE_OFN18_n4568), 
	.A1(FE_OFN1627_acc_fft_data_in_0_), 
	.A0(n8473));
   AO22XLTS U1942 (.Y(n6164), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[14] ), 
	.B0(FE_OFN11_n4568), 
	.A1(FE_OFN1547_acc_fft_data_in_14_), 
	.A0(n8476));
   AO22XLTS U1946 (.Y(n6168), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[10] ), 
	.B0(FE_OFN13_n4568), 
	.A1(FE_OFN1567_acc_fft_data_in_10_), 
	.A0(n8475));
   AO22XLTS U1941 (.Y(n6163), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[15] ), 
	.B0(FE_OFN11_n4568), 
	.A1(FE_OFN1540_acc_fft_data_in_15_), 
	.A0(n8476));
   AO22XLTS U1947 (.Y(n6169), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[9] ), 
	.B0(FE_OFN14_n4568), 
	.A1(FE_OFN1572_acc_fft_data_in_9_), 
	.A0(n8475));
   AO22XLTS U1952 (.Y(n6174), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[4] ), 
	.B0(FE_OFN19_n4568), 
	.A1(FE_OFN1602_acc_fft_data_in_4_), 
	.A0(n8474));
   AO22XLTS U1944 (.Y(n6166), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[12] ), 
	.B0(FE_OFN10_n4568), 
	.A1(FE_OFN1557_acc_fft_data_in_12_), 
	.A0(n8476));
   AO22XLTS U1943 (.Y(n6165), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[13] ), 
	.B0(FE_OFN11_n4568), 
	.A1(FE_OFN1552_acc_fft_data_in_13_), 
	.A0(n8476));
   AO22XLTS U1954 (.Y(n6176), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[2] ), 
	.B0(FE_OFN21_n4568), 
	.A1(FE_OFN1613_acc_fft_data_in_2_), 
	.A0(n8473));
   AO22XLTS U1955 (.Y(n6177), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[1] ), 
	.B0(FE_OFN21_n4568), 
	.A1(FE_OFN1618_acc_fft_data_in_1_), 
	.A0(n8473));
   AO22XLTS U1945 (.Y(n6167), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[11] ), 
	.B0(FE_OFN14_n4568), 
	.A1(FE_OFN1562_acc_fft_data_in_11_), 
	.A0(n8475));
   OAI211XLTS U1063 (.Y(n4168), 
	.C0(n9474), 
	.B0(\fifo_to_fir/hang[3] ), 
	.A1(n4170), 
	.A0(n8790));
   OAI211XLTS U919 (.Y(n3993), 
	.C0(n9478), 
	.B0(\fifo_to_fft/hang[3] ), 
	.A1(n3995), 
	.A0(n8811));
   AO22XLTS U1953 (.Y(n6175), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[3] ), 
	.B0(FE_OFN20_n4568), 
	.A1(FE_OFN1606_acc_fft_data_in_3_), 
	.A0(n8473));
   AO22XLTS U1948 (.Y(n6170), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[8] ), 
	.B0(FE_OFN14_n4568), 
	.A1(FE_OFN1576_acc_fft_data_in_8_), 
	.A0(n8475));
   AO22XLTS U1951 (.Y(n6173), 
	.B1(\fifo_from_fft/fifo_cell2/sr_out[5] ), 
	.B0(FE_OFN19_n4568), 
	.A1(FE_OFN1595_acc_fft_data_in_5_), 
	.A0(n8474));
   CLKINVX1TS U615 (.Y(n5351), 
	.A(n3719));
   CLKINVX1TS U623 (.Y(n5355), 
	.A(n3726));
   CLKINVX1TS U625 (.Y(n5356), 
	.A(n3727));
   CLKINVX1TS U617 (.Y(n5352), 
	.A(n3723));
   CLKINVX1TS U627 (.Y(n5357), 
	.A(n3728));
   CLKINVX1TS U629 (.Y(n5358), 
	.A(n3729));
   CLKINVX1TS U621 (.Y(n5354), 
	.A(n3725));
   CLKINVX1TS U619 (.Y(n5353), 
	.A(n3724));
   CLKINVX1TS U647 (.Y(n5367), 
	.A(n3738));
   CLKINVX1TS U649 (.Y(n5368), 
	.A(n3739));
   CLKINVX1TS U651 (.Y(n5369), 
	.A(n3740));
   CLKINVX1TS U653 (.Y(n5370), 
	.A(n3741));
   CLKINVX1TS U655 (.Y(n5371), 
	.A(n3742));
   AOI22X1TS U467 (.Y(n3624), 
	.B1(\router/addr_calc/fft_write_calc/counter/N72 ), 
	.B0(FE_OFN954_n3619), 
	.A1(FE_OFN971_n3618), 
	.A0(n7377));
   CLKINVX1TS U657 (.Y(n5372), 
	.A(n3743));
   CLKINVX1TS U659 (.Y(n5373), 
	.A(n3744));
   CLKINVX1TS U661 (.Y(n5374), 
	.A(n3745));
   NAND2XLTS U346 (.Y(\router/addr_calc/fir_write_calc/counter/N189 ), 
	.B(n3551), 
	.A(n9417));
   AOI22X1TS U317 (.Y(n3536), 
	.B1(\router/addr_calc/fir_write_calc/counter/N72 ), 
	.B0(FE_OFN894_n3531), 
	.A1(FE_OFN900_n3530), 
	.A0(n7135));
   NAND2XLTS U443 (.Y(\router/addr_calc/fir_read_calc/counter/N178 ), 
	.B(n3606), 
	.A(n9407));
   NAND2XLTS U421 (.Y(\router/addr_calc/fir_read_calc/counter/N189 ), 
	.B(n3595), 
	.A(n9410));
   AOI22X1TS U392 (.Y(n3580), 
	.B1(\router/addr_calc/fir_read_calc/counter/N72 ), 
	.B0(FE_OFN917_n3575), 
	.A1(FE_OFN928_n3574), 
	.A0(n7263));
   AOI22X1TS U542 (.Y(n3668), 
	.B1(\router/addr_calc/fft_read_calc/counter/N72 ), 
	.B0(FE_OFN868_n3663), 
	.A1(FE_OFN880_n3662), 
	.A0(n7501));
   NAND2XLTS U425 (.Y(\router/addr_calc/fir_read_calc/counter/N187 ), 
	.B(n3597), 
	.A(n9413));
   NAND2XLTS U350 (.Y(\router/addr_calc/fir_write_calc/counter/N187 ), 
	.B(n3553), 
	.A(n9417));
   AOI22X1TS U242 (.Y(n3492), 
	.B1(\router/addr_calc/iir_write_calc/counter/N72 ), 
	.B0(FE_OFN930_n3487), 
	.A1(FE_OFN943_n3486), 
	.A0(n7180));
   OAI21XLTS U2554 (.Y(n4749), 
	.B0(FE_OFN653_n4747), 
	.A1(n4752), 
	.A0(n7589));
   AOI22X1TS U465 (.Y(n3623), 
	.B1(\router/addr_calc/fft_write_calc/counter/N73 ), 
	.B0(FE_OFN954_n3619), 
	.A1(FE_OFN972_n3618), 
	.A0(\router/addr_calc/fft_write_calc/count[27] ));
   AOI22X1TS U240 (.Y(n3491), 
	.B1(\router/addr_calc/iir_write_calc/counter/N73 ), 
	.B0(FE_OFN933_n3487), 
	.A1(FE_OFN943_n3486), 
	.A0(FE_OFN1439_router_addr_calc_iir_write_calc_count_27_));
   AOI22X1TS U390 (.Y(n3579), 
	.B1(\router/addr_calc/fir_read_calc/counter/N73 ), 
	.B0(FE_OFN918_n3575), 
	.A1(FE_OFN928_n3574), 
	.A0(FE_OFN1239_router_addr_calc_fir_read_calc_count_27_));
   AOI22X1TS U315 (.Y(n3535), 
	.B1(\router/addr_calc/fir_write_calc/counter/N73 ), 
	.B0(FE_OFN894_n3531), 
	.A1(FE_OFN900_n3530), 
	.A0(\router/addr_calc/fir_write_calc/count[27] ));
   AOI22X1TS U540 (.Y(n3667), 
	.B1(\router/addr_calc/fft_read_calc/counter/N73 ), 
	.B0(FE_OFN868_n3663), 
	.A1(FE_OFN879_n3662), 
	.A0(FE_OFN1237_router_addr_calc_fft_read_calc_count_27_));
   NAND3XLTS U2678 (.Y(n4649), 
	.C(n4820), 
	.B(n4650), 
	.A(FE_OFN654_n4747));
   OAI21X1TS U1923 (.Y(n4563), 
	.B0(FE_OFN313_n4561), 
	.A1(n4566), 
	.A0(n7514));
   AOI21X1TS U2552 (.Y(n6674), 
	.B0(FE_OFN828_n7619), 
	.A1(n4749), 
	.A0(\fifo_from_fir/fifo_cell3/controller/valid_read ));
   OAI21XLTS U2553 (.Y(n6675), 
	.B0(n4749), 
	.A1(n4751), 
	.A0(\fifo_from_fir/fifo_cell3/data_out/N35 ));
   AOI22X1TS U463 (.Y(n3622), 
	.B1(\router/addr_calc/fft_write_calc/counter/N74 ), 
	.B0(FE_OFN952_n3619), 
	.A1(FE_OFN972_n3618), 
	.A0(n7372));
   AOI22X1TS U388 (.Y(n3578), 
	.B1(\router/addr_calc/fir_read_calc/counter/N74 ), 
	.B0(FE_OFN917_n3575), 
	.A1(FE_OFN928_n3574), 
	.A0(n7258));
   AOI22X1TS U538 (.Y(n3666), 
	.B1(\router/addr_calc/fft_read_calc/counter/N74 ), 
	.B0(FE_OFN870_n3663), 
	.A1(FE_OFN879_n3662), 
	.A0(n7496));
   AOI22X1TS U238 (.Y(n3490), 
	.B1(\router/addr_calc/iir_write_calc/counter/N74 ), 
	.B0(FE_OFN933_n3487), 
	.A1(FE_OFN941_n3486), 
	.A0(n7186));
   AOI22X1TS U313 (.Y(n3534), 
	.B1(\router/addr_calc/fir_write_calc/counter/N74 ), 
	.B0(FE_OFN893_n3531), 
	.A1(FE_OFN900_n3530), 
	.A0(n7129));
   AO22XLTS U2521 (.Y(n6644), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[29] ), 
	.B0(FE_OFN367_n4748), 
	.A1(FE_OFN1643_acc_fir_data_in_29_), 
	.A0(FE_OFN657_n4747));
   AO22XLTS U2522 (.Y(n6645), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[28] ), 
	.B0(FE_OFN367_n4748), 
	.A1(FE_OFN1648_acc_fir_data_in_28_), 
	.A0(FE_OFN657_n4747));
   AO22XLTS U2519 (.Y(n6642), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[31] ), 
	.B0(FE_OFN367_n4748), 
	.A1(FE_OFN1630_acc_fir_data_in_31_), 
	.A0(FE_OFN657_n4747));
   AO22XLTS U2520 (.Y(n6643), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[30] ), 
	.B0(FE_OFN367_n4748), 
	.A1(FE_OFN1635_acc_fir_data_in_30_), 
	.A0(FE_OFN655_n4747));
   AO22XLTS U2536 (.Y(n6659), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[14] ), 
	.B0(FE_OFN368_n4748), 
	.A1(FE_OFN1730_acc_fir_data_in_14_), 
	.A0(FE_OFN663_n4747));
   AO22XLTS U2537 (.Y(n6660), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[13] ), 
	.B0(FE_OFN363_n4748), 
	.A1(FE_OFN1733_acc_fir_data_in_13_), 
	.A0(FE_OFN661_n4747));
   AO22XLTS U2538 (.Y(n6661), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[12] ), 
	.B0(FE_OFN368_n4748), 
	.A1(FE_OFN1739_acc_fir_data_in_12_), 
	.A0(FE_OFN663_n4747));
   AOI21X1TS U1921 (.Y(n6145), 
	.B0(FE_OFN818_n7619), 
	.A1(n4563), 
	.A0(\fifo_from_fft/fifo_cell3/controller/valid_read ));
   NAND3XLTS U2047 (.Y(n4463), 
	.C(n4634), 
	.B(n4464), 
	.A(n4561));
   AO22XLTS U2535 (.Y(n6658), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[15] ), 
	.B0(FE_OFN368_n4748), 
	.A1(FE_OFN1723_acc_fir_data_in_15_), 
	.A0(FE_OFN663_n4747));
   OAI211XLTS U2679 (.Y(n4819), 
	.C0(n9466), 
	.B0(\fifo_from_fir/hang[2] ), 
	.A1(n4821), 
	.A0(n8876));
   OAI21XLTS U1922 (.Y(n6146), 
	.B0(n4563), 
	.A1(n4565), 
	.A0(\fifo_from_fft/fifo_cell3/data_out/N35 ));
   AOI22X1TS U536 (.Y(n3665), 
	.B1(\router/addr_calc/fft_read_calc/counter/N75 ), 
	.B0(FE_OFN870_n3663), 
	.A1(FE_OFN878_n3662), 
	.A0(FE_OFN1234_n7492));
   AOI22X1TS U386 (.Y(n3577), 
	.B1(\router/addr_calc/fir_read_calc/counter/N75 ), 
	.B0(FE_OFN918_n3575), 
	.A1(FE_OFN929_n3574), 
	.A0(FE_OFN1235_n7254));
   AOI22X1TS U311 (.Y(n3533), 
	.B1(\router/addr_calc/fir_write_calc/counter/N75 ), 
	.B0(FE_OFN894_n3531), 
	.A1(FE_OFN899_n3530), 
	.A0(n7124));
   AOI22X1TS U461 (.Y(n3621), 
	.B1(\router/addr_calc/fft_write_calc/counter/N75 ), 
	.B0(FE_OFN952_n3619), 
	.A1(FE_OFN972_n3618), 
	.A0(\router/addr_calc/fft_write_calc/count[29] ));
   AOI22X1TS U236 (.Y(n3489), 
	.B1(\router/addr_calc/iir_write_calc/counter/N75 ), 
	.B0(FE_OFN933_n3487), 
	.A1(FE_OFN941_n3486), 
	.A0(n7192));
   AO22XLTS U1896 (.Y(n6121), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[23] ), 
	.B0(FE_OFN23_n4562), 
	.A1(FE_OFN1494_acc_fft_data_in_23_), 
	.A0(FE_OFN316_n4561));
   OAI21XLTS U1011 (.Y(n5552), 
	.B0(n4110), 
	.A1(n4109), 
	.A0(\fifo_to_fir/fifo_cell5/data_out/N35 ));
   AO22XLTS U1898 (.Y(n6123), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[21] ), 
	.B0(FE_OFN27_n4562), 
	.A1(FE_OFN1508_acc_fft_data_in_21_), 
	.A0(FE_OFN319_n4561));
   OAI21XLTS U867 (.Y(n5500), 
	.B0(n3935), 
	.A1(n3934), 
	.A0(\fifo_to_fft/fifo_cell5/data_out/N35 ));
   OAI211XLTS U2048 (.Y(n4633), 
	.C0(n9470), 
	.B0(\fifo_from_fft/hang[2] ), 
	.A1(n4635), 
	.A0(n8843));
   AO22XLTS U1888 (.Y(n6113), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[31] ), 
	.B0(FE_OFN27_n4562), 
	.A1(FE_OFN1456_acc_fft_data_in_31_), 
	.A0(FE_OFN317_n4561));
   AO22XLTS U1897 (.Y(n6122), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[22] ), 
	.B0(FE_OFN29_n4562), 
	.A1(FE_OFN1503_acc_fft_data_in_22_), 
	.A0(FE_OFN319_n4561));
   AO22XLTS U2550 (.Y(n6673), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[0] ), 
	.B0(FE_OFN359_n4748), 
	.A1(FE_OFN1814_acc_fir_data_in_0_), 
	.A0(FE_OFN656_n4747));
   AO22XLTS U1889 (.Y(n6114), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[30] ), 
	.B0(FE_OFN28_n4562), 
	.A1(FE_OFN1462_acc_fft_data_in_30_), 
	.A0(FE_OFN321_n4561));
   AOI21X1TS U869 (.Y(n5501), 
	.B0(FE_OFN826_n7619), 
	.A1(n3935), 
	.A0(\fifo_to_fft/fifo_cell5/controller/valid_read ));
   AO22XLTS U2549 (.Y(n6672), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[1] ), 
	.B0(FE_OFN359_n4748), 
	.A1(FE_OFN1804_acc_fir_data_in_1_), 
	.A0(FE_OFN656_n4747));
   AO22XLTS U1899 (.Y(n6124), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[20] ), 
	.B0(FE_OFN29_n4562), 
	.A1(FE_OFN1514_acc_fft_data_in_20_), 
	.A0(FE_OFN322_n4561));
   AO22XLTS U2527 (.Y(n6650), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[23] ), 
	.B0(FE_OFN360_n4748), 
	.A1(FE_OFN1673_acc_fir_data_in_23_), 
	.A0(FE_OFN659_n4747));
   AO22XLTS U2548 (.Y(n6671), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[2] ), 
	.B0(FE_OFN359_n4748), 
	.A1(FE_OFN1797_acc_fir_data_in_2_), 
	.A0(FE_OFN656_n4747));
   AO22XLTS U2547 (.Y(n6670), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[3] ), 
	.B0(n4748), 
	.A1(FE_OFN1792_acc_fir_data_in_3_), 
	.A0(FE_OFN658_n4747));
   AO22XLTS U2546 (.Y(n6669), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[4] ), 
	.B0(FE_OFN362_n4748), 
	.A1(FE_OFN1784_acc_fir_data_in_4_), 
	.A0(FE_OFN654_n4747));
   AO22XLTS U2545 (.Y(n6668), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[5] ), 
	.B0(FE_OFN364_n4748), 
	.A1(FE_OFN1780_acc_fir_data_in_5_), 
	.A0(n4747));
   AO22XLTS U1890 (.Y(n6115), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[29] ), 
	.B0(FE_OFN26_n4562), 
	.A1(FE_OFN1467_acc_fft_data_in_29_), 
	.A0(FE_OFN318_n4561));
   AO22XLTS U2544 (.Y(n6667), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[6] ), 
	.B0(FE_OFN364_n4748), 
	.A1(FE_OFN1769_acc_fir_data_in_6_), 
	.A0(FE_OFN657_n4747));
   AO22XLTS U2543 (.Y(n6666), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[7] ), 
	.B0(FE_OFN362_n4748), 
	.A1(FE_OFN1768_acc_fir_data_in_7_), 
	.A0(FE_OFN654_n4747));
   AO22XLTS U2542 (.Y(n6665), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[8] ), 
	.B0(FE_OFN366_n4748), 
	.A1(FE_OFN1761_acc_fir_data_in_8_), 
	.A0(FE_OFN662_n4747));
   AO22XLTS U2541 (.Y(n6664), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[9] ), 
	.B0(FE_OFN366_n4748), 
	.A1(FE_OFN1754_acc_fir_data_in_9_), 
	.A0(FE_OFN662_n4747));
   AO22XLTS U1891 (.Y(n6116), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[28] ), 
	.B0(FE_OFN27_n4562), 
	.A1(FE_OFN1471_acc_fft_data_in_28_), 
	.A0(FE_OFN318_n4561));
   AO22XLTS U2540 (.Y(n6663), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[10] ), 
	.B0(FE_OFN366_n4748), 
	.A1(FE_OFN1747_acc_fir_data_in_10_), 
	.A0(FE_OFN662_n4747));
   AO22XLTS U2539 (.Y(n6662), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[11] ), 
	.B0(FE_OFN363_n4748), 
	.A1(FE_OFN1745_acc_fir_data_in_11_), 
	.A0(FE_OFN661_n4747));
   NAND3XLTS U916 (.Y(n3860), 
	.C(n3991), 
	.B(n3861), 
	.A(n7315));
   AO22XLTS U2530 (.Y(n6653), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[20] ), 
	.B0(FE_OFN360_n4748), 
	.A1(FE_OFN1694_acc_fir_data_in_20_), 
	.A0(FE_OFN659_n4747));
   NAND3XLTS U1060 (.Y(n4035), 
	.C(n4166), 
	.B(n4036), 
	.A(n7424));
   AO22XLTS U2523 (.Y(n6646), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[27] ), 
	.B0(FE_OFN365_n4748), 
	.A1(FE_OFN1653_acc_fir_data_in_27_), 
	.A0(FE_OFN655_n4747));
   AO22XLTS U2524 (.Y(n6647), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[26] ), 
	.B0(FE_OFN365_n4748), 
	.A1(FE_OFN1818_acc_fir_data_in_26_), 
	.A0(FE_OFN655_n4747));
   AO22XLTS U2533 (.Y(n6656), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[17] ), 
	.B0(FE_OFN361_n4748), 
	.A1(FE_OFN1708_acc_fir_data_in_17_), 
	.A0(FE_OFN660_n4747));
   AO22XLTS U2525 (.Y(n6648), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[25] ), 
	.B0(FE_OFN365_n4748), 
	.A1(FE_OFN1661_acc_fir_data_in_25_), 
	.A0(FE_OFN652_n4747));
   AO22XLTS U2529 (.Y(n6652), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[21] ), 
	.B0(FE_OFN360_n4748), 
	.A1(FE_OFN1683_acc_fir_data_in_21_), 
	.A0(FE_OFN660_n4747));
   AO22XLTS U2531 (.Y(n6654), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[19] ), 
	.B0(n4748), 
	.A1(FE_OFN1701_acc_fir_data_in_19_), 
	.A0(FE_OFN659_n4747));
   AO22XLTS U2534 (.Y(n6657), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[16] ), 
	.B0(FE_OFN361_n4748), 
	.A1(FE_OFN1716_acc_fir_data_in_16_), 
	.A0(FE_OFN660_n4747));
   AO22XLTS U2526 (.Y(n6649), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[24] ), 
	.B0(FE_OFN365_n4748), 
	.A1(FE_OFN1666_acc_fir_data_in_24_), 
	.A0(FE_OFN652_n4747));
   AO22XLTS U2528 (.Y(n6651), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[22] ), 
	.B0(FE_OFN368_n4748), 
	.A1(FE_OFN1682_acc_fir_data_in_22_), 
	.A0(FE_OFN663_n4747));
   AO22XLTS U2532 (.Y(n6655), 
	.B1(\fifo_from_fir/fifo_cell3/sr_out[18] ), 
	.B0(FE_OFN363_n4748), 
	.A1(FE_OFN1703_acc_fir_data_in_18_), 
	.A0(FE_OFN661_n4747));
   AOI22X1TS U309 (.Y(n3532), 
	.B1(\router/addr_calc/fir_write_calc/counter/N76 ), 
	.B0(FE_OFN897_n3531), 
	.A1(n3530), 
	.A0(FE_OFN1231_router_addr_calc_fir_write_calc_count_30_));
   AOI22X1TS U234 (.Y(n3488), 
	.B1(\router/addr_calc/iir_write_calc/counter/N76 ), 
	.B0(FE_OFN933_n3487), 
	.A1(FE_OFN941_n3486), 
	.A0(\router/addr_calc/iir_write_calc/count[30] ));
   AOI22X1TS U384 (.Y(n3576), 
	.B1(\router/addr_calc/fir_read_calc/counter/N76 ), 
	.B0(FE_OFN918_n3575), 
	.A1(FE_OFN929_n3574), 
	.A0(\router/addr_calc/fir_read_calc/count[30] ));
   AOI22X1TS U534 (.Y(n3664), 
	.B1(\router/addr_calc/fft_read_calc/counter/N76 ), 
	.B0(FE_OFN873_n3663), 
	.A1(FE_OFN879_n3662), 
	.A0(\router/addr_calc/fft_read_calc/count[30] ));
   AOI22X1TS U459 (.Y(n3620), 
	.B1(\router/addr_calc/fft_write_calc/counter/N76 ), 
	.B0(FE_OFN960_n3619), 
	.A1(FE_OFN963_n3618), 
	.A0(FE_OFN1232_n7368));
   AO22XLTS U1914 (.Y(n6139), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[5] ), 
	.B0(FE_OFN26_n4562), 
	.A1(FE_OFN1591_acc_fft_data_in_5_), 
	.A0(FE_OFN317_n4561));
   AO22XLTS U1908 (.Y(n6133), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[11] ), 
	.B0(FE_OFN31_n4562), 
	.A1(FE_OFN1563_acc_fft_data_in_11_), 
	.A0(FE_OFN322_n4561));
   AO22XLTS U1915 (.Y(n6140), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[4] ), 
	.B0(FE_OFN22_n4562), 
	.A1(FE_OFN1600_acc_fft_data_in_4_), 
	.A0(FE_OFN314_n4561));
   AO22XLTS U1906 (.Y(n6131), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[13] ), 
	.B0(FE_OFN30_n4562), 
	.A1(FE_OFN1549_acc_fft_data_in_13_), 
	.A0(FE_OFN323_n4561));
   AO22XLTS U1901 (.Y(n6126), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[18] ), 
	.B0(FE_OFN23_n4562), 
	.A1(FE_OFN1520_acc_fft_data_in_18_), 
	.A0(FE_OFN316_n4561));
   AO22XLTS U1893 (.Y(n6118), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[26] ), 
	.B0(FE_OFN28_n4562), 
	.A1(FE_OFN1479_acc_fft_data_in_26_), 
	.A0(FE_OFN321_n4561));
   AO22XLTS U1910 (.Y(n6135), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[9] ), 
	.B0(FE_OFN31_n4562), 
	.A1(FE_OFN1570_acc_fft_data_in_9_), 
	.A0(FE_OFN322_n4561));
   AO22XLTS U1905 (.Y(n6130), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[14] ), 
	.B0(FE_OFN32_n4562), 
	.A1(FE_OFN1544_acc_fft_data_in_14_), 
	.A0(FE_OFN324_n4561));
   OAI211XLTS U1061 (.Y(n4165), 
	.C0(n9472), 
	.B0(\fifo_to_fir/hang[4] ), 
	.A1(n4167), 
	.A0(n8790));
   AO22XLTS U1904 (.Y(n6129), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[15] ), 
	.B0(FE_OFN30_n4562), 
	.A1(FE_OFN1542_acc_fft_data_in_15_), 
	.A0(FE_OFN323_n4561));
   AO22XLTS U1900 (.Y(n6125), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[19] ), 
	.B0(n4562), 
	.A1(FE_OFN1517_acc_fft_data_in_19_), 
	.A0(FE_OFN313_n4561));
   AO22XLTS U1909 (.Y(n6134), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[10] ), 
	.B0(FE_OFN29_n4562), 
	.A1(FE_OFN1567_acc_fft_data_in_10_), 
	.A0(FE_OFN319_n4561));
   AO22XLTS U1911 (.Y(n6136), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[8] ), 
	.B0(FE_OFN31_n4562), 
	.A1(FE_OFN1576_acc_fft_data_in_8_), 
	.A0(FE_OFN323_n4561));
   AO22XLTS U1916 (.Y(n6141), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[3] ), 
	.B0(FE_OFN28_n4562), 
	.A1(FE_OFN1603_acc_fft_data_in_3_), 
	.A0(FE_OFN321_n4561));
   AO22XLTS U1913 (.Y(n6138), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[6] ), 
	.B0(FE_OFN23_n4562), 
	.A1(FE_OFN1586_acc_fft_data_in_6_), 
	.A0(FE_OFN316_n4561));
   AO22XLTS U1895 (.Y(n6120), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[24] ), 
	.B0(FE_OFN25_n4562), 
	.A1(FE_OFN1489_acc_fft_data_in_24_), 
	.A0(FE_OFN320_n4561));
   AO22XLTS U1917 (.Y(n6142), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[2] ), 
	.B0(FE_OFN25_n4562), 
	.A1(FE_OFN1609_acc_fft_data_in_2_), 
	.A0(FE_OFN320_n4561));
   AO22XLTS U1892 (.Y(n6117), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[27] ), 
	.B0(FE_OFN24_n4562), 
	.A1(FE_OFN1474_acc_fft_data_in_27_), 
	.A0(FE_OFN315_n4561));
   AO22XLTS U1907 (.Y(n6132), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[12] ), 
	.B0(FE_OFN32_n4562), 
	.A1(FE_OFN1555_acc_fft_data_in_12_), 
	.A0(FE_OFN324_n4561));
   AO22XLTS U1918 (.Y(n6143), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[1] ), 
	.B0(FE_OFN24_n4562), 
	.A1(FE_OFN1616_acc_fft_data_in_1_), 
	.A0(FE_OFN315_n4561));
   AO22XLTS U1912 (.Y(n6137), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[7] ), 
	.B0(FE_OFN22_n4562), 
	.A1(FE_OFN1583_acc_fft_data_in_7_), 
	.A0(FE_OFN315_n4561));
   OAI211XLTS U917 (.Y(n3990), 
	.C0(n9476), 
	.B0(\fifo_to_fft/hang[4] ), 
	.A1(n3992), 
	.A0(n8811));
   AO22XLTS U1903 (.Y(n6128), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[16] ), 
	.B0(FE_OFN32_n4562), 
	.A1(FE_OFN1533_acc_fft_data_in_16_), 
	.A0(FE_OFN324_n4561));
   AO22XLTS U1919 (.Y(n6144), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[0] ), 
	.B0(FE_OFN28_n4562), 
	.A1(FE_OFN1627_acc_fft_data_in_0_), 
	.A0(FE_OFN321_n4561));
   AO22XLTS U1894 (.Y(n6119), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[25] ), 
	.B0(FE_OFN25_n4562), 
	.A1(FE_OFN1486_acc_fft_data_in_25_), 
	.A0(FE_OFN320_n4561));
   AO22XLTS U1902 (.Y(n6127), 
	.B1(\fifo_from_fft/fifo_cell3/sr_out[17] ), 
	.B0(FE_OFN32_n4562), 
	.A1(FE_OFN1529_acc_fft_data_in_17_), 
	.A0(FE_OFN324_n4561));
   AOI22X1TS U382 (.Y(n3573), 
	.B1(\router/addr_calc/fir_read_calc/counter/N77 ), 
	.B0(FE_OFN918_n3575), 
	.A1(FE_OFN929_n3574), 
	.A0(n7249));
   AOI22X1TS U457 (.Y(n3617), 
	.B1(\router/addr_calc/fft_write_calc/counter/N77 ), 
	.B0(FE_OFN952_n3619), 
	.A1(FE_OFN972_n3618), 
	.A0(\router/addr_calc/fft_write_calc/count[31] ));
   AOI22X1TS U307 (.Y(n3529), 
	.B1(\router/addr_calc/fir_write_calc/counter/N77 ), 
	.B0(FE_OFN897_n3531), 
	.A1(FE_OFN898_n3530), 
	.A0(n7118));
   AOI22X1TS U532 (.Y(n3661), 
	.B1(\router/addr_calc/fft_read_calc/counter/N77 ), 
	.B0(FE_OFN875_n3663), 
	.A1(FE_OFN877_n3662), 
	.A0(n7487));
   OAI21X1TS U2517 (.Y(n4743), 
	.B0(FE_OFN642_n4741), 
	.A1(n4746), 
	.A0(n7584));
   NAND2XLTS U306 (.Y(\router/addr_calc/fir_write_calc/counter/N209 ), 
	.B(n3529), 
	.A(n9407));
   AO22XLTS U2509 (.Y(n6635), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[4] ), 
	.B0(FE_OFN632_n4742), 
	.A1(FE_OFN1787_acc_fir_data_in_4_), 
	.A0(FE_OFN640_n4741));
   AOI21X1TS U2515 (.Y(n6640), 
	.B0(FE_OFN829_n7619), 
	.A1(n4743), 
	.A0(\fifo_from_fir/fifo_cell4/controller/valid_read ));
   NAND3XLTS U2676 (.Y(n4651), 
	.C(n4817), 
	.B(n4652), 
	.A(FE_OFN642_n4741));
   NAND3XLTS U914 (.Y(n3862), 
	.C(n3988), 
	.B(n3863), 
	.A(n3932));
   OAI21XLTS U2516 (.Y(n6641), 
	.B0(n4743), 
	.A1(n4745), 
	.A0(\fifo_from_fir/fifo_cell4/data_out/N35 ));
   NAND3XLTS U1058 (.Y(n4037), 
	.C(n4163), 
	.B(n4038), 
	.A(n4107));
   OAI21X1TS U1886 (.Y(n4557), 
	.B0(FE_OFN301_n4555), 
	.A1(n4560), 
	.A0(n7509));
   AOI21X1TS U864 (.Y(n5498), 
	.B0(FE_OFN834_n7619), 
	.A1(n3930), 
	.A0(\fifo_to_fft/fifo_cell6/controller/valid_read ));
   AOI21X1TS U1008 (.Y(n5550), 
	.B0(FE_OFN811_n7619), 
	.A1(n4105), 
	.A0(\fifo_to_fir/fifo_cell6/controller/valid_read ));
   OAI21XLTS U1885 (.Y(n6112), 
	.B0(n4557), 
	.A1(n4559), 
	.A0(\fifo_from_fft/fifo_cell4/data_out/N35 ));
   AO22XLTS U2506 (.Y(n6632), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[7] ), 
	.B0(FE_OFN632_n4742), 
	.A1(FE_OFN1768_acc_fir_data_in_7_), 
	.A0(FE_OFN640_n4741));
   OAI211XLTS U915 (.Y(n3987), 
	.C0(n9477), 
	.B0(\fifo_to_fft/hang[5] ), 
	.A1(n3989), 
	.A0(n8811));
   OAI21XLTS U1006 (.Y(n5549), 
	.B0(n4105), 
	.A1(n4104), 
	.A0(\fifo_to_fir/fifo_cell6/data_out/N35 ));
   AO22XLTS U2507 (.Y(n6633), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[6] ), 
	.B0(FE_OFN638_n4742), 
	.A1(FE_OFN1771_acc_fir_data_in_6_), 
	.A0(FE_OFN645_n4741));
   OAI211XLTS U1059 (.Y(n4162), 
	.C0(n9474), 
	.B0(\fifo_to_fir/hang[5] ), 
	.A1(n4164), 
	.A0(n8790));
   AOI21X1TS U1884 (.Y(n6111), 
	.B0(FE_OFN825_n7619), 
	.A1(n4557), 
	.A0(\fifo_from_fft/fifo_cell4/controller/valid_read ));
   AO22XLTS U2508 (.Y(n6634), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[5] ), 
	.B0(FE_OFN632_n4742), 
	.A1(FE_OFN1779_acc_fir_data_in_5_), 
	.A0(n4741));
   OAI211XLTS U2677 (.Y(n4816), 
	.C0(n9466), 
	.B0(\fifo_from_fir/hang[3] ), 
	.A1(n4818), 
	.A0(n8876));
   NAND3XLTS U2045 (.Y(n4465), 
	.C(n4631), 
	.B(n4466), 
	.A(n4555));
   OAI21XLTS U862 (.Y(n5497), 
	.B0(n3930), 
	.A1(n3929), 
	.A0(\fifo_to_fft/fifo_cell6/data_out/N35 ));
   AO22XLTS U1878 (.Y(n6106), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[4] ), 
	.B0(n4556), 
	.A1(FE_OFN1599_acc_fft_data_in_4_), 
	.A0(FE_OFN301_n4555));
   AO22XLTS U2497 (.Y(n6623), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[16] ), 
	.B0(FE_OFN630_n4742), 
	.A1(FE_OFN1717_acc_fir_data_in_16_), 
	.A0(FE_OFN647_n4741));
   AO22XLTS U2495 (.Y(n6621), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[18] ), 
	.B0(FE_OFN634_n4742), 
	.A1(FE_OFN1706_acc_fir_data_in_18_), 
	.A0(FE_OFN649_n4741));
   AO22XLTS U2494 (.Y(n6620), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[19] ), 
	.B0(n4742), 
	.A1(FE_OFN1699_acc_fir_data_in_19_), 
	.A0(FE_OFN647_n4741));
   AO22XLTS U2496 (.Y(n6622), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[17] ), 
	.B0(FE_OFN630_n4742), 
	.A1(FE_OFN1711_acc_fir_data_in_17_), 
	.A0(FE_OFN647_n4741));
   AO22XLTS U2493 (.Y(n6619), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[20] ), 
	.B0(FE_OFN630_n4742), 
	.A1(FE_OFN1690_acc_fir_data_in_20_), 
	.A0(FE_OFN648_n4741));
   AO22XLTS U2513 (.Y(n6639), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[0] ), 
	.B0(n4742), 
	.A1(FE_OFN1816_acc_fir_data_in_0_), 
	.A0(FE_OFN646_n4741));
   AO22XLTS U2492 (.Y(n6618), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[21] ), 
	.B0(FE_OFN634_n4742), 
	.A1(FE_OFN1684_acc_fir_data_in_21_), 
	.A0(FE_OFN648_n4741));
   AO22XLTS U2512 (.Y(n6638), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[1] ), 
	.B0(FE_OFN631_n4742), 
	.A1(FE_OFN1803_acc_fir_data_in_1_), 
	.A0(FE_OFN644_n4741));
   AO22XLTS U2510 (.Y(n6636), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[3] ), 
	.B0(FE_OFN631_n4742), 
	.A1(FE_OFN1794_acc_fir_data_in_3_), 
	.A0(FE_OFN644_n4741));
   AO22XLTS U2511 (.Y(n6637), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[2] ), 
	.B0(FE_OFN631_n4742), 
	.A1(FE_OFN1801_acc_fir_data_in_2_), 
	.A0(FE_OFN644_n4741));
   AO22XLTS U2490 (.Y(n6616), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[23] ), 
	.B0(FE_OFN634_n4742), 
	.A1(FE_OFN1677_acc_fir_data_in_23_), 
	.A0(FE_OFN648_n4741));
   AO22XLTS U2491 (.Y(n6617), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[22] ), 
	.B0(FE_OFN639_n4742), 
	.A1(FE_OFN1682_acc_fir_data_in_22_), 
	.A0(FE_OFN651_n4741));
   OAI21XLTS U860 (.Y(n3925), 
	.B0(n3927), 
	.A1(n3923), 
	.A0(n7301));
   AO22XLTS U1875 (.Y(n6103), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[7] ), 
	.B0(FE_OFN299_n4556), 
	.A1(FE_OFN1581_acc_fft_data_in_7_), 
	.A0(FE_OFN308_n4555));
   AO22XLTS U1876 (.Y(n6104), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[6] ), 
	.B0(FE_OFN291_n4556), 
	.A1(FE_OFN1587_acc_fft_data_in_6_), 
	.A0(FE_OFN303_n4555));
   OAI21XLTS U1004 (.Y(n4100), 
	.B0(n4102), 
	.A1(n4098), 
	.A0(n7410));
   OAI211XLTS U2046 (.Y(n4630), 
	.C0(n9470), 
	.B0(\fifo_from_fft/hang[3] ), 
	.A1(n4632), 
	.A0(n8843));
   AO22XLTS U1877 (.Y(n6105), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[5] ), 
	.B0(FE_OFN294_n4556), 
	.A1(FE_OFN1593_acc_fft_data_in_5_), 
	.A0(FE_OFN305_n4555));
   NAND3XLTS U1056 (.Y(n4039), 
	.C(n4160), 
	.B(n4040), 
	.A(n4102));
   AO22XLTS U1881 (.Y(n6109), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[1] ), 
	.B0(FE_OFN294_n4556), 
	.A1(FE_OFN1615_acc_fft_data_in_1_), 
	.A0(FE_OFN305_n4555));
   OAI21XLTS U857 (.Y(n5494), 
	.B0(n3925), 
	.A1(n3924), 
	.A0(\fifo_to_fft/fifo_cell7/data_out/N35 ));
   AO22XLTS U1879 (.Y(n6107), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[3] ), 
	.B0(FE_OFN300_n4556), 
	.A1(FE_OFN1603_acc_fft_data_in_3_), 
	.A0(FE_OFN309_n4555));
   AO22XLTS U1880 (.Y(n6108), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[2] ), 
	.B0(FE_OFN299_n4556), 
	.A1(FE_OFN1608_acc_fft_data_in_2_), 
	.A0(FE_OFN308_n4555));
   AO22XLTS U1882 (.Y(n6110), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[0] ), 
	.B0(FE_OFN300_n4556), 
	.A1(FE_OFN1627_acc_fft_data_in_0_), 
	.A0(FE_OFN309_n4555));
   AO22XLTS U2499 (.Y(n6625), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[14] ), 
	.B0(FE_OFN639_n4742), 
	.A1(FE_OFN1730_acc_fir_data_in_14_), 
	.A0(FE_OFN651_n4741));
   AO22XLTS U2500 (.Y(n6626), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[13] ), 
	.B0(FE_OFN633_n4742), 
	.A1(FE_OFN1735_acc_fir_data_in_13_), 
	.A0(FE_OFN649_n4741));
   AO22XLTS U2501 (.Y(n6627), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[12] ), 
	.B0(FE_OFN639_n4742), 
	.A1(FE_OFN1739_acc_fir_data_in_12_), 
	.A0(FE_OFN651_n4741));
   OAI21XLTS U1001 (.Y(n5546), 
	.B0(n4100), 
	.A1(n4099), 
	.A0(\fifo_to_fir/fifo_cell7/data_out/N35 ));
   AO22XLTS U2502 (.Y(n6628), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[11] ), 
	.B0(FE_OFN633_n4742), 
	.A1(FE_OFN1744_acc_fir_data_in_11_), 
	.A0(FE_OFN649_n4741));
   AO22XLTS U2503 (.Y(n6629), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[10] ), 
	.B0(FE_OFN636_n4742), 
	.A1(FE_OFN1749_acc_fir_data_in_10_), 
	.A0(FE_OFN650_n4741));
   AO22XLTS U2504 (.Y(n6630), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[9] ), 
	.B0(FE_OFN636_n4742), 
	.A1(FE_OFN1754_acc_fir_data_in_9_), 
	.A0(FE_OFN650_n4741));
   NAND3XLTS U912 (.Y(n3864), 
	.C(n3985), 
	.B(n3865), 
	.A(n3927));
   AO22XLTS U1861 (.Y(n6089), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[21] ), 
	.B0(FE_OFN295_n4556), 
	.A1(FE_OFN1508_acc_fft_data_in_21_), 
	.A0(FE_OFN306_n4555));
   AOI21X1TS U1003 (.Y(n5547), 
	.B0(FE_OFN800_n7619), 
	.A1(n4100), 
	.A0(\fifo_to_fir/fifo_cell7/controller/valid_read ));
   AO22XLTS U1862 (.Y(n6090), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[20] ), 
	.B0(FE_OFN293_n4556), 
	.A1(FE_OFN1510_acc_fft_data_in_20_), 
	.A0(FE_OFN310_n4555));
   AO22XLTS U1864 (.Y(n6092), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[18] ), 
	.B0(n4556), 
	.A1(FE_OFN1523_acc_fft_data_in_18_), 
	.A0(FE_OFN302_n4555));
   AO22XLTS U2484 (.Y(n6610), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[29] ), 
	.B0(FE_OFN638_n4742), 
	.A1(FE_OFN1645_acc_fir_data_in_29_), 
	.A0(FE_OFN645_n4741));
   AO22XLTS U1863 (.Y(n6091), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[19] ), 
	.B0(n4556), 
	.A1(FE_OFN1518_acc_fft_data_in_19_), 
	.A0(FE_OFN302_n4555));
   AO22XLTS U1859 (.Y(n6087), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[23] ), 
	.B0(FE_OFN291_n4556), 
	.A1(FE_OFN1494_acc_fft_data_in_23_), 
	.A0(FE_OFN303_n4555));
   AO22XLTS U2486 (.Y(n6612), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[27] ), 
	.B0(FE_OFN635_n4742), 
	.A1(FE_OFN1655_acc_fir_data_in_27_), 
	.A0(FE_OFN643_n4741));
   AO22XLTS U2482 (.Y(n6608), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[31] ), 
	.B0(FE_OFN638_n4742), 
	.A1(FE_OFN1631_acc_fir_data_in_31_), 
	.A0(FE_OFN645_n4741));
   AOI21X1TS U859 (.Y(n5495), 
	.B0(FE_OFN797_n7619), 
	.A1(n3925), 
	.A0(\fifo_to_fft/fifo_cell7/controller/valid_read ));
   AO22XLTS U2489 (.Y(n6615), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[24] ), 
	.B0(FE_OFN637_n4742), 
	.A1(FE_OFN1670_acc_fir_data_in_24_), 
	.A0(FE_OFN641_n4741));
   AO22XLTS U2488 (.Y(n6614), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[25] ), 
	.B0(FE_OFN637_n4742), 
	.A1(FE_OFN1665_acc_fir_data_in_25_), 
	.A0(FE_OFN643_n4741));
   AO22XLTS U2487 (.Y(n6613), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[26] ), 
	.B0(FE_OFN637_n4742), 
	.A1(FE_OFN1658_acc_fir_data_in_26_), 
	.A0(FE_OFN641_n4741));
   AO22XLTS U2483 (.Y(n6609), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[30] ), 
	.B0(FE_OFN635_n4742), 
	.A1(FE_OFN1637_acc_fir_data_in_30_), 
	.A0(FE_OFN643_n4741));
   AO22XLTS U2505 (.Y(n6631), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[8] ), 
	.B0(FE_OFN636_n4742), 
	.A1(FE_OFN1761_acc_fir_data_in_8_), 
	.A0(FE_OFN650_n4741));
   AO22XLTS U1860 (.Y(n6088), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[22] ), 
	.B0(FE_OFN295_n4556), 
	.A1(FE_OFN1503_acc_fft_data_in_22_), 
	.A0(FE_OFN306_n4555));
   AO22XLTS U1865 (.Y(n6093), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[17] ), 
	.B0(FE_OFN297_n4556), 
	.A1(FE_OFN1528_acc_fft_data_in_17_), 
	.A0(FE_OFN312_n4555));
   AO22XLTS U1866 (.Y(n6094), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[16] ), 
	.B0(FE_OFN297_n4556), 
	.A1(FE_OFN1533_acc_fft_data_in_16_), 
	.A0(FE_OFN312_n4555));
   AO22XLTS U2485 (.Y(n6611), 
	.B1(\fifo_from_fir/fifo_cell4/sr_out[28] ), 
	.B0(FE_OFN638_n4742), 
	.A1(FE_OFN1650_acc_fir_data_in_28_), 
	.A0(FE_OFN645_n4741));
   AO22XLTS U1852 (.Y(n6080), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[30] ), 
	.B0(FE_OFN300_n4556), 
	.A1(FE_OFN1462_acc_fft_data_in_30_), 
	.A0(FE_OFN309_n4555));
   AO22XLTS U1853 (.Y(n6081), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[29] ), 
	.B0(FE_OFN300_n4556), 
	.A1(FE_OFN1467_acc_fft_data_in_29_), 
	.A0(FE_OFN309_n4555));
   AO22XLTS U1854 (.Y(n6082), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[28] ), 
	.B0(FE_OFN295_n4556), 
	.A1(FE_OFN1471_acc_fft_data_in_28_), 
	.A0(FE_OFN304_n4555));
   OAI211XLTS U913 (.Y(n3984), 
	.C0(n9478), 
	.B0(\fifo_to_fft/hang[6] ), 
	.A1(n3986), 
	.A0(n8810));
   AO22XLTS U1851 (.Y(n6079), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[31] ), 
	.B0(FE_OFN295_n4556), 
	.A1(FE_OFN1454_acc_fft_data_in_31_), 
	.A0(FE_OFN304_n4555));
   AO22XLTS U1857 (.Y(n6085), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[25] ), 
	.B0(FE_OFN299_n4556), 
	.A1(FE_OFN1483_acc_fft_data_in_25_), 
	.A0(FE_OFN308_n4555));
   AO22XLTS U1855 (.Y(n6083), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[27] ), 
	.B0(FE_OFN298_n4556), 
	.A1(FE_OFN1473_acc_fft_data_in_27_), 
	.A0(FE_OFN307_n4555));
   AO22XLTS U1872 (.Y(n6100), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[10] ), 
	.B0(FE_OFN292_n4556), 
	.A1(FE_OFN1567_acc_fft_data_in_10_), 
	.A0(FE_OFN306_n4555));
   AO22XLTS U1858 (.Y(n6086), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[24] ), 
	.B0(FE_OFN299_n4556), 
	.A1(FE_OFN1488_acc_fft_data_in_24_), 
	.A0(FE_OFN308_n4555));
   AO22XLTS U1870 (.Y(n6098), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[12] ), 
	.B0(FE_OFN297_n4556), 
	.A1(FE_OFN1555_acc_fft_data_in_12_), 
	.A0(FE_OFN312_n4555));
   AO22XLTS U1873 (.Y(n6101), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[9] ), 
	.B0(FE_OFN296_n4556), 
	.A1(FE_OFN1570_acc_fft_data_in_9_), 
	.A0(FE_OFN310_n4555));
   OAI211XLTS U1057 (.Y(n4159), 
	.C0(n9474), 
	.B0(\fifo_to_fir/hang[6] ), 
	.A1(n4161), 
	.A0(n8789));
   AO22XLTS U1868 (.Y(n6096), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[14] ), 
	.B0(FE_OFN297_n4556), 
	.A1(FE_OFN1543_acc_fft_data_in_14_), 
	.A0(FE_OFN312_n4555));
   AO22XLTS U1871 (.Y(n6099), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[11] ), 
	.B0(FE_OFN296_n4556), 
	.A1(FE_OFN1563_acc_fft_data_in_11_), 
	.A0(FE_OFN310_n4555));
   AO22XLTS U1869 (.Y(n6097), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[13] ), 
	.B0(FE_OFN296_n4556), 
	.A1(FE_OFN1548_acc_fft_data_in_13_), 
	.A0(FE_OFN311_n4555));
   AO22XLTS U1874 (.Y(n6102), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[8] ), 
	.B0(FE_OFN296_n4556), 
	.A1(FE_OFN1575_acc_fft_data_in_8_), 
	.A0(FE_OFN311_n4555));
   AO22XLTS U1856 (.Y(n6084), 
	.B1(\fifo_from_fft/fifo_cell4/sr_out[26] ), 
	.B0(FE_OFN298_n4556), 
	.A1(FE_OFN1479_acc_fft_data_in_26_), 
	.A0(FE_OFN307_n4555));
   OAI21X1TS U2480 (.Y(n4737), 
	.B0(FE_OFN618_n4735), 
	.A1(n4740), 
	.A0(n7579));
   OAI21XLTS U1849 (.Y(n4551), 
	.B0(n4549), 
	.A1(n4554), 
	.A0(n7504));
   AOI21X1TS U2478 (.Y(n6606), 
	.B0(FE_OFN829_n7619), 
	.A1(n4737), 
	.A0(\fifo_from_fir/fifo_cell5/controller/valid_read ));
   NAND3XLTS U2674 (.Y(n4653), 
	.C(n4814), 
	.B(n4654), 
	.A(FE_OFN618_n4735));
   OAI21XLTS U2479 (.Y(n6607), 
	.B0(n4737), 
	.A1(n4739), 
	.A0(\fifo_from_fir/fifo_cell5/data_out/N35 ));
   OAI21XLTS U1848 (.Y(n6078), 
	.B0(n4551), 
	.A1(n4553), 
	.A0(\fifo_from_fft/fifo_cell5/data_out/N35 ));
   AO22XLTS U2463 (.Y(n6592), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[13] ), 
	.B0(FE_OFN374_n4736), 
	.A1(FE_OFN1734_acc_fir_data_in_13_), 
	.A0(FE_OFN627_n4735));
   NAND3XLTS U2043 (.Y(n4467), 
	.C(n4628), 
	.B(n4468), 
	.A(n4549));
   AO22XLTS U2446 (.Y(n6575), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[30] ), 
	.B0(FE_OFN375_n4736), 
	.A1(FE_OFN1636_acc_fir_data_in_30_), 
	.A0(FE_OFN624_n4735));
   AO22XLTS U2464 (.Y(n6593), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[12] ), 
	.B0(FE_OFN378_n4736), 
	.A1(FE_OFN1739_acc_fir_data_in_12_), 
	.A0(FE_OFN629_n4735));
   AO22XLTS U2461 (.Y(n6590), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[15] ), 
	.B0(FE_OFN378_n4736), 
	.A1(FE_OFN1723_acc_fir_data_in_15_), 
	.A0(FE_OFN629_n4735));
   AO22XLTS U2448 (.Y(n6577), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[28] ), 
	.B0(FE_OFN375_n4736), 
	.A1(FE_OFN1649_acc_fir_data_in_28_), 
	.A0(FE_OFN623_n4735));
   AO22XLTS U2447 (.Y(n6576), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[29] ), 
	.B0(FE_OFN375_n4736), 
	.A1(FE_OFN1644_acc_fir_data_in_29_), 
	.A0(FE_OFN623_n4735));
   AO22XLTS U2462 (.Y(n6591), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[14] ), 
	.B0(FE_OFN378_n4736), 
	.A1(FE_OFN1730_acc_fir_data_in_14_), 
	.A0(FE_OFN629_n4735));
   AO22XLTS U2445 (.Y(n6574), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[31] ), 
	.B0(FE_OFN373_n4736), 
	.A1(FE_OFN1630_acc_fir_data_in_31_), 
	.A0(FE_OFN623_n4735));
   AOI21X1TS U1847 (.Y(n6077), 
	.B0(FE_OFN832_n7619), 
	.A1(n4551), 
	.A0(\fifo_from_fft/fifo_cell5/controller/valid_read ));
   OAI211XLTS U2675 (.Y(n4813), 
	.C0(n9466), 
	.B0(\fifo_from_fir/hang[4] ), 
	.A1(n4815), 
	.A0(n8876));
   AO22XLTS U2476 (.Y(n6605), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[0] ), 
	.B0(FE_OFN370_n4736), 
	.A1(FE_OFN1813_acc_fir_data_in_0_), 
	.A0(FE_OFN619_n4735));
   AO22XLTS U2471 (.Y(n6600), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[5] ), 
	.B0(FE_OFN372_n4736), 
	.A1(FE_OFN1780_acc_fir_data_in_5_), 
	.A0(n4735));
   AO22XLTS U2472 (.Y(n6601), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[4] ), 
	.B0(FE_OFN372_n4736), 
	.A1(FE_OFN1787_acc_fir_data_in_4_), 
	.A0(n4735));
   AO22XLTS U2473 (.Y(n6602), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[3] ), 
	.B0(FE_OFN370_n4736), 
	.A1(FE_OFN1793_acc_fir_data_in_3_), 
	.A0(FE_OFN621_n4735));
   AO22XLTS U2468 (.Y(n6597), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[8] ), 
	.B0(FE_OFN376_n4736), 
	.A1(FE_OFN1761_acc_fir_data_in_8_), 
	.A0(FE_OFN628_n4735));
   AO22XLTS U1814 (.Y(n6045), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[31] ), 
	.B0(FE_OFN36_n4550), 
	.A1(FE_OFN1454_acc_fft_data_in_31_), 
	.A0(FE_OFN285_n4549));
   AO22XLTS U2466 (.Y(n6595), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[10] ), 
	.B0(FE_OFN376_n4736), 
	.A1(FE_OFN1749_acc_fir_data_in_10_), 
	.A0(FE_OFN628_n4735));
   AO22XLTS U2465 (.Y(n6594), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[11] ), 
	.B0(FE_OFN374_n4736), 
	.A1(FE_OFN1744_acc_fir_data_in_11_), 
	.A0(FE_OFN627_n4735));
   AO22XLTS U2470 (.Y(n6599), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[6] ), 
	.B0(FE_OFN373_n4736), 
	.A1(FE_OFN1771_acc_fir_data_in_6_), 
	.A0(FE_OFN620_n4735));
   AO22XLTS U2475 (.Y(n6604), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[1] ), 
	.B0(FE_OFN370_n4736), 
	.A1(FE_OFN1806_acc_fir_data_in_1_), 
	.A0(FE_OFN621_n4735));
   AO22XLTS U1815 (.Y(n6046), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[30] ), 
	.B0(FE_OFN35_n4550), 
	.A1(FE_OFN1459_acc_fft_data_in_30_), 
	.A0(FE_OFN286_n4549));
   AO22XLTS U2474 (.Y(n6603), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[2] ), 
	.B0(FE_OFN372_n4736), 
	.A1(FE_OFN1800_acc_fir_data_in_2_), 
	.A0(FE_OFN619_n4735));
   AO22XLTS U2460 (.Y(n6589), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[16] ), 
	.B0(FE_OFN371_n4736), 
	.A1(FE_OFN1718_acc_fir_data_in_16_), 
	.A0(FE_OFN625_n4735));
   AO22XLTS U2467 (.Y(n6596), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[9] ), 
	.B0(FE_OFN376_n4736), 
	.A1(FE_OFN1754_acc_fir_data_in_9_), 
	.A0(FE_OFN628_n4735));
   AO22XLTS U2459 (.Y(n6588), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[17] ), 
	.B0(FE_OFN369_n4736), 
	.A1(FE_OFN1710_acc_fir_data_in_17_), 
	.A0(FE_OFN622_n4735));
   AO22XLTS U1830 (.Y(n6061), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[15] ), 
	.B0(FE_OFN39_n4550), 
	.A1(FE_OFN1539_acc_fft_data_in_15_), 
	.A0(FE_OFN282_n4549));
   OAI211XLTS U2044 (.Y(n4627), 
	.C0(n9468), 
	.B0(\fifo_from_fft/hang[4] ), 
	.A1(n4629), 
	.A0(n8843));
   AO22XLTS U2458 (.Y(n6587), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[18] ), 
	.B0(FE_OFN374_n4736), 
	.A1(FE_OFN1705_acc_fir_data_in_18_), 
	.A0(FE_OFN627_n4735));
   AO22XLTS U2457 (.Y(n6586), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[19] ), 
	.B0(FE_OFN369_n4736), 
	.A1(FE_OFN1701_acc_fir_data_in_19_), 
	.A0(FE_OFN622_n4735));
   AO22XLTS U2456 (.Y(n6585), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[20] ), 
	.B0(FE_OFN369_n4736), 
	.A1(FE_OFN1694_acc_fir_data_in_20_), 
	.A0(FE_OFN622_n4735));
   AO22XLTS U2455 (.Y(n6584), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[21] ), 
	.B0(FE_OFN371_n4736), 
	.A1(FE_OFN1683_acc_fir_data_in_21_), 
	.A0(FE_OFN625_n4735));
   AO22XLTS U2469 (.Y(n6598), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[7] ), 
	.B0(FE_OFN373_n4736), 
	.A1(FE_OFN1765_acc_fir_data_in_7_), 
	.A0(FE_OFN620_n4735));
   AO22XLTS U2454 (.Y(n6583), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[22] ), 
	.B0(FE_OFN378_n4736), 
	.A1(FE_OFN1682_acc_fir_data_in_22_), 
	.A0(FE_OFN629_n4735));
   AO22XLTS U2453 (.Y(n6582), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[23] ), 
	.B0(FE_OFN371_n4736), 
	.A1(FE_OFN1672_acc_fir_data_in_23_), 
	.A0(FE_OFN625_n4735));
   AO22XLTS U1816 (.Y(n6047), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[29] ), 
	.B0(FE_OFN36_n4550), 
	.A1(FE_OFN1465_acc_fft_data_in_29_), 
	.A0(FE_OFN286_n4549));
   AO22XLTS U1817 (.Y(n6048), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[28] ), 
	.B0(FE_OFN36_n4550), 
	.A1(FE_OFN1820_acc_fft_data_in_28_), 
	.A0(FE_OFN285_n4549));
   AO22XLTS U2452 (.Y(n6581), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[24] ), 
	.B0(FE_OFN377_n4736), 
	.A1(FE_OFN1668_acc_fir_data_in_24_), 
	.A0(FE_OFN626_n4735));
   AO22XLTS U1831 (.Y(n6062), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[14] ), 
	.B0(FE_OFN40_n4550), 
	.A1(FE_OFN1544_acc_fft_data_in_14_), 
	.A0(FE_OFN282_n4549));
   AO22XLTS U2451 (.Y(n6580), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[25] ), 
	.B0(FE_OFN377_n4736), 
	.A1(FE_OFN1662_acc_fir_data_in_25_), 
	.A0(FE_OFN626_n4735));
   AO22XLTS U2450 (.Y(n6579), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[26] ), 
	.B0(FE_OFN377_n4736), 
	.A1(FE_OFN1660_acc_fir_data_in_26_), 
	.A0(FE_OFN624_n4735));
   AO22XLTS U1833 (.Y(n6064), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[12] ), 
	.B0(FE_OFN41_n4550), 
	.A1(FE_OFN1555_acc_fft_data_in_12_), 
	.A0(FE_OFN280_n4549));
   AO22XLTS U1832 (.Y(n6063), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[13] ), 
	.B0(FE_OFN39_n4550), 
	.A1(FE_OFN1550_acc_fft_data_in_13_), 
	.A0(FE_OFN282_n4549));
   AO22XLTS U2449 (.Y(n6578), 
	.B1(\fifo_from_fir/fifo_cell5/sr_out[27] ), 
	.B0(FE_OFN377_n4736), 
	.A1(FE_OFN1654_acc_fir_data_in_27_), 
	.A0(FE_OFN624_n4735));
   AO22XLTS U1823 (.Y(n6054), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[22] ), 
	.B0(FE_OFN37_n4550), 
	.A1(FE_OFN1499_acc_fft_data_in_22_), 
	.A0(FE_OFN284_n4549));
   AO22XLTS U1845 (.Y(n6076), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[0] ), 
	.B0(FE_OFN35_n4550), 
	.A1(FE_OFN1627_acc_fft_data_in_0_), 
	.A0(FE_OFN286_n4549));
   AO22XLTS U1829 (.Y(n6060), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[16] ), 
	.B0(FE_OFN41_n4550), 
	.A1(FE_OFN1534_acc_fft_data_in_16_), 
	.A0(FE_OFN280_n4549));
   AO22XLTS U1824 (.Y(n6055), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[21] ), 
	.B0(FE_OFN37_n4550), 
	.A1(FE_OFN1506_acc_fft_data_in_21_), 
	.A0(FE_OFN285_n4549));
   AO22XLTS U1836 (.Y(n6067), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[9] ), 
	.B0(FE_OFN38_n4550), 
	.A1(FE_OFN1570_acc_fft_data_in_9_), 
	.A0(FE_OFN283_n4549));
   AO22XLTS U1844 (.Y(n6075), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[1] ), 
	.B0(FE_OFN34_n4550), 
	.A1(FE_OFN1617_acc_fft_data_in_1_), 
	.A0(FE_OFN288_n4549));
   AO22XLTS U1839 (.Y(n6070), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[6] ), 
	.B0(FE_OFN42_n4550), 
	.A1(FE_OFN1585_acc_fft_data_in_6_), 
	.A0(FE_OFN281_n4549));
   AO22XLTS U1826 (.Y(n6057), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[19] ), 
	.B0(FE_OFN42_n4550), 
	.A1(FE_OFN1516_acc_fft_data_in_19_), 
	.A0(FE_OFN279_n4549));
   AO22XLTS U1837 (.Y(n6068), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[8] ), 
	.B0(FE_OFN38_n4550), 
	.A1(FE_OFN1575_acc_fft_data_in_8_), 
	.A0(FE_OFN283_n4549));
   AO22XLTS U1842 (.Y(n6073), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[3] ), 
	.B0(FE_OFN35_n4550), 
	.A1(FE_OFN1606_acc_fft_data_in_3_), 
	.A0(FE_OFN287_n4549));
   AO22XLTS U1835 (.Y(n6066), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[10] ), 
	.B0(FE_OFN38_n4550), 
	.A1(FE_OFN1566_acc_fft_data_in_10_), 
	.A0(FE_OFN284_n4549));
   NAND3XLTS U910 (.Y(n3866), 
	.C(n3982), 
	.B(n3867), 
	.A(n7295));
   AO22XLTS U1818 (.Y(n6049), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[27] ), 
	.B0(FE_OFN34_n4550), 
	.A1(FE_OFN1475_acc_fft_data_in_27_), 
	.A0(FE_OFN287_n4549));
   AO22XLTS U1838 (.Y(n6069), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[7] ), 
	.B0(n4550), 
	.A1(FE_OFN1581_acc_fft_data_in_7_), 
	.A0(FE_OFN290_n4549));
   AO22XLTS U1820 (.Y(n6051), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[25] ), 
	.B0(FE_OFN33_n4550), 
	.A1(FE_OFN1486_acc_fft_data_in_25_), 
	.A0(FE_OFN289_n4549));
   AO22XLTS U1841 (.Y(n6072), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[4] ), 
	.B0(n4550), 
	.A1(FE_OFN1600_acc_fft_data_in_4_), 
	.A0(FE_OFN290_n4549));
   OAI21XLTS U996 (.Y(n5543), 
	.B0(n4095), 
	.A1(n4094), 
	.A0(\fifo_to_fir/fifo_cell8/data_out/N35 ));
   AO22XLTS U1843 (.Y(n6074), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[2] ), 
	.B0(FE_OFN33_n4550), 
	.A1(FE_OFN1610_acc_fft_data_in_2_), 
	.A0(FE_OFN288_n4549));
   AO22XLTS U1840 (.Y(n6071), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[5] ), 
	.B0(FE_OFN42_n4550), 
	.A1(FE_OFN1591_acc_fft_data_in_5_), 
	.A0(FE_OFN281_n4549));
   AO22XLTS U1821 (.Y(n6052), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[24] ), 
	.B0(FE_OFN33_n4550), 
	.A1(FE_OFN1489_acc_fft_data_in_24_), 
	.A0(FE_OFN288_n4549));
   AO22XLTS U1828 (.Y(n6059), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[17] ), 
	.B0(FE_OFN41_n4550), 
	.A1(FE_OFN1528_acc_fft_data_in_17_), 
	.A0(FE_OFN280_n4549));
   AO22XLTS U1834 (.Y(n6065), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[11] ), 
	.B0(FE_OFN39_n4550), 
	.A1(FE_OFN1563_acc_fft_data_in_11_), 
	.A0(FE_OFN283_n4549));
   AO22XLTS U1819 (.Y(n6050), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[26] ), 
	.B0(FE_OFN34_n4550), 
	.A1(FE_OFN1480_acc_fft_data_in_26_), 
	.A0(FE_OFN287_n4549));
   AO22XLTS U1827 (.Y(n6058), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[18] ), 
	.B0(FE_OFN40_n4550), 
	.A1(FE_OFN1526_acc_fft_data_in_18_), 
	.A0(FE_OFN281_n4549));
   AO22XLTS U1825 (.Y(n6056), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[20] ), 
	.B0(FE_OFN37_n4550), 
	.A1(FE_OFN1514_acc_fft_data_in_20_), 
	.A0(FE_OFN284_n4549));
   OAI21XLTS U852 (.Y(n5491), 
	.B0(n3920), 
	.A1(n3919), 
	.A0(\fifo_to_fft/fifo_cell8/data_out/N35 ));
   AO22XLTS U1822 (.Y(n6053), 
	.B1(\fifo_from_fft/fifo_cell5/sr_out[23] ), 
	.B0(FE_OFN42_n4550), 
	.A1(FE_OFN1493_acc_fft_data_in_23_), 
	.A0(FE_OFN281_n4549));
   NAND3XLTS U1054 (.Y(n4041), 
	.C(n4157), 
	.B(n4042), 
	.A(n7404));
   OAI211XLTS U1055 (.Y(n4156), 
	.C0(n9475), 
	.B0(\fifo_to_fir/hang[7] ), 
	.A1(n4158), 
	.A0(n8789));
   OAI211XLTS U911 (.Y(n3981), 
	.C0(n9479), 
	.B0(\fifo_to_fft/hang[7] ), 
	.A1(n3983), 
	.A0(n8810));
   OAI21XLTS U2443 (.Y(n4731), 
	.B0(n4729), 
	.A1(n4734), 
	.A0(n7574));
   OAI21XLTS U1812 (.Y(n4545), 
	.B0(n4543), 
	.A1(n4548), 
	.A0(n7499));
   NAND3XLTS U2672 (.Y(n4655), 
	.C(n4811), 
	.B(n4656), 
	.A(n4729));
   AO22XLTS U2418 (.Y(n6550), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[21] ), 
	.B0(FE_OFN381_n4730), 
	.A1(FE_OFN1684_acc_fir_data_in_21_), 
	.A0(FE_OFN614_n4729));
   AOI21X1TS U2441 (.Y(n6572), 
	.B0(FE_OFN822_n7619), 
	.A1(n4731), 
	.A0(\fifo_from_fir/fifo_cell6/controller/valid_read ));
   OAI21XLTS U2442 (.Y(n6573), 
	.B0(n4731), 
	.A1(n4733), 
	.A0(\fifo_from_fir/fifo_cell6/data_out/N35 ));
   AO22XLTS U2417 (.Y(n6549), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[22] ), 
	.B0(FE_OFN389_n4730), 
	.A1(FE_OFN1681_acc_fir_data_in_22_), 
	.A0(FE_OFN617_n4729));
   AO22XLTS U2419 (.Y(n6551), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[20] ), 
	.B0(FE_OFN381_n4730), 
	.A1(FE_OFN1690_acc_fir_data_in_20_), 
	.A0(FE_OFN610_n4729));
   AO22XLTS U2416 (.Y(n6548), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[23] ), 
	.B0(FE_OFN381_n4730), 
	.A1(FE_OFN1677_acc_fir_data_in_23_), 
	.A0(FE_OFN610_n4729));
   AOI21X1TS U1810 (.Y(n6043), 
	.B0(FE_OFN832_n7619), 
	.A1(n4545), 
	.A0(\fifo_from_fft/fifo_cell6/controller/valid_read ));
   AO22XLTS U2408 (.Y(n6540), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[31] ), 
	.B0(FE_OFN388_n4730), 
	.A1(FE_OFN1629_acc_fir_data_in_31_), 
	.A0(FE_OFN613_n4729));
   AO22XLTS U1786 (.Y(n6020), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[22] ), 
	.B0(FE_OFN265_n4544), 
	.A1(FE_OFN1499_acc_fft_data_in_22_), 
	.A0(FE_OFN275_n4543));
   OAI21XLTS U1811 (.Y(n6044), 
	.B0(n4545), 
	.A1(n4547), 
	.A0(\fifo_from_fft/fifo_cell6/data_out/N35 ));
   AO22XLTS U1787 (.Y(n6021), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[21] ), 
	.B0(FE_OFN264_n4544), 
	.A1(FE_OFN1506_acc_fft_data_in_21_), 
	.A0(FE_OFN275_n4543));
   AO22XLTS U2410 (.Y(n6542), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[29] ), 
	.B0(FE_OFN388_n4730), 
	.A1(FE_OFN1640_acc_fir_data_in_29_), 
	.A0(FE_OFN613_n4729));
   AO22XLTS U2409 (.Y(n6541), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[30] ), 
	.B0(FE_OFN388_n4730), 
	.A1(FE_OFN1634_acc_fir_data_in_30_), 
	.A0(FE_OFN613_n4729));
   OAI211XLTS U2673 (.Y(n4810), 
	.C0(n9467), 
	.B0(\fifo_from_fir/hang[5] ), 
	.A1(n4812), 
	.A0(n8876));
   NAND3XLTS U2041 (.Y(n4469), 
	.C(n4625), 
	.B(n4470), 
	.A(n4543));
   NAND3XLTS U908 (.Y(n3868), 
	.C(n3979), 
	.B(n3869), 
	.A(n7285));
   AO22XLTS U1779 (.Y(n6013), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[29] ), 
	.B0(FE_OFN263_n4544), 
	.A1(FE_OFN1463_acc_fft_data_in_29_), 
	.A0(FE_OFN277_n4543));
   AO22XLTS U1785 (.Y(n6019), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[23] ), 
	.B0(FE_OFN265_n4544), 
	.A1(FE_OFN1495_acc_fft_data_in_23_), 
	.A0(FE_OFN271_n4543));
   AO22XLTS U1788 (.Y(n6022), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[20] ), 
	.B0(FE_OFN265_n4544), 
	.A1(FE_OFN1513_acc_fft_data_in_20_), 
	.A0(FE_OFN271_n4543));
   AO22XLTS U1778 (.Y(n6012), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[30] ), 
	.B0(FE_OFN263_n4544), 
	.A1(FE_OFN1459_acc_fft_data_in_30_), 
	.A0(FE_OFN277_n4543));
   OAI21XLTS U847 (.Y(n5488), 
	.B0(n3915), 
	.A1(n3914), 
	.A0(\fifo_to_fft/fifo_cell9/data_out/N35 ));
   AO22XLTS U2422 (.Y(n6554), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[17] ), 
	.B0(FE_OFN383_n4730), 
	.A1(FE_OFN1708_acc_fir_data_in_17_), 
	.A0(FE_OFN614_n4729));
   AO22XLTS U2411 (.Y(n6543), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[28] ), 
	.B0(FE_OFN388_n4730), 
	.A1(FE_OFN1647_acc_fir_data_in_28_), 
	.A0(FE_OFN613_n4729));
   AO22XLTS U2423 (.Y(n6555), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[16] ), 
	.B0(FE_OFN383_n4730), 
	.A1(FE_OFN1715_acc_fir_data_in_16_), 
	.A0(FE_OFN614_n4729));
   OAI211XLTS U2042 (.Y(n4624), 
	.C0(n9470), 
	.B0(\fifo_from_fft/hang[5] ), 
	.A1(n4626), 
	.A0(n8843));
   AO22XLTS U2421 (.Y(n6553), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[18] ), 
	.B0(FE_OFN384_n4730), 
	.A1(FE_OFN1704_acc_fir_data_in_18_), 
	.A0(FE_OFN615_n4729));
   OAI21XLTS U991 (.Y(n5540), 
	.B0(n4090), 
	.A1(n4089), 
	.A0(\fifo_to_fir/fifo_cell9/data_out/N35 ));
   AO22XLTS U1777 (.Y(n6011), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[31] ), 
	.B0(FE_OFN264_n4544), 
	.A1(FE_OFN1457_acc_fft_data_in_31_), 
	.A0(FE_OFN277_n4543));
   AO22XLTS U2420 (.Y(n6552), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[19] ), 
	.B0(FE_OFN379_n4730), 
	.A1(FE_OFN1701_acc_fir_data_in_19_), 
	.A0(FE_OFN610_n4729));
   NAND3XLTS U1052 (.Y(n4043), 
	.C(n4154), 
	.B(n4044), 
	.A(n7394));
   AO22XLTS U1790 (.Y(n6024), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[18] ), 
	.B0(FE_OFN257_n4544), 
	.A1(FE_OFN1526_acc_fft_data_in_18_), 
	.A0(FE_OFN267_n4543));
   AO22XLTS U1791 (.Y(n6025), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[17] ), 
	.B0(FE_OFN257_n4544), 
	.A1(FE_OFN1527_acc_fft_data_in_17_), 
	.A0(FE_OFN266_n4543));
   AO22XLTS U1792 (.Y(n6026), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[16] ), 
	.B0(FE_OFN257_n4544), 
	.A1(FE_OFN1534_acc_fft_data_in_16_), 
	.A0(FE_OFN266_n4543));
   AO22XLTS U1780 (.Y(n6014), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[28] ), 
	.B0(FE_OFN264_n4544), 
	.A1(FE_OFN1468_acc_fft_data_in_28_), 
	.A0(FE_OFN277_n4543));
   OAI211XLTS U1053 (.Y(n4153), 
	.C0(n9475), 
	.B0(\fifo_to_fir/hang[8] ), 
	.A1(n4155), 
	.A0(n8789));
   AO22XLTS U1789 (.Y(n6023), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[19] ), 
	.B0(n4544), 
	.A1(FE_OFN1517_acc_fft_data_in_19_), 
	.A0(FE_OFN267_n4543));
   OAI211XLTS U909 (.Y(n3978), 
	.C0(n9478), 
	.B0(\fifo_to_fft/hang[8] ), 
	.A1(n3980), 
	.A0(n8810));
   AO22XLTS U2439 (.Y(n6571), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[0] ), 
	.B0(FE_OFN380_n4730), 
	.A1(FE_OFN1816_acc_fir_data_in_0_), 
	.A0(FE_OFN608_n4729));
   AO22XLTS U2426 (.Y(n6558), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[13] ), 
	.B0(FE_OFN384_n4730), 
	.A1(FE_OFN1732_acc_fir_data_in_13_), 
	.A0(FE_OFN615_n4729));
   AO22XLTS U2425 (.Y(n6557), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[14] ), 
	.B0(FE_OFN389_n4730), 
	.A1(FE_OFN1725_acc_fir_data_in_14_), 
	.A0(FE_OFN617_n4729));
   AO22XLTS U2438 (.Y(n6570), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[1] ), 
	.B0(n4730), 
	.A1(FE_OFN1806_acc_fir_data_in_1_), 
	.A0(FE_OFN606_n4729));
   AO22XLTS U2437 (.Y(n6569), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[2] ), 
	.B0(FE_OFN380_n4730), 
	.A1(FE_OFN1801_acc_fir_data_in_2_), 
	.A0(FE_OFN609_n4729));
   AO22XLTS U2436 (.Y(n6568), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[3] ), 
	.B0(n4730), 
	.A1(FE_OFN1793_acc_fir_data_in_3_), 
	.A0(FE_OFN606_n4729));
   AO22XLTS U2435 (.Y(n6567), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[4] ), 
	.B0(FE_OFN382_n4730), 
	.A1(FE_OFN1787_acc_fir_data_in_4_), 
	.A0(FE_OFN607_n4729));
   AO22XLTS U2434 (.Y(n6566), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[5] ), 
	.B0(FE_OFN385_n4730), 
	.A1(FE_OFN1780_acc_fir_data_in_5_), 
	.A0(FE_OFN607_n4729));
   AO22XLTS U2433 (.Y(n6565), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[6] ), 
	.B0(FE_OFN382_n4730), 
	.A1(FE_OFN1769_acc_fir_data_in_6_), 
	.A0(FE_OFN609_n4729));
   AO22XLTS U2432 (.Y(n6564), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[7] ), 
	.B0(FE_OFN382_n4730), 
	.A1(FE_OFN1763_acc_fir_data_in_7_), 
	.A0(FE_OFN609_n4729));
   AO22XLTS U2431 (.Y(n6563), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[8] ), 
	.B0(FE_OFN387_n4730), 
	.A1(FE_OFN1759_acc_fir_data_in_8_), 
	.A0(FE_OFN616_n4729));
   AO22XLTS U2430 (.Y(n6562), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[9] ), 
	.B0(FE_OFN387_n4730), 
	.A1(FE_OFN1752_acc_fir_data_in_9_), 
	.A0(FE_OFN616_n4729));
   AO22XLTS U2429 (.Y(n6561), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[10] ), 
	.B0(FE_OFN387_n4730), 
	.A1(FE_OFN1749_acc_fir_data_in_10_), 
	.A0(FE_OFN616_n4729));
   AO22XLTS U2428 (.Y(n6560), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[11] ), 
	.B0(FE_OFN384_n4730), 
	.A1(FE_OFN1745_acc_fir_data_in_11_), 
	.A0(FE_OFN615_n4729));
   AO22XLTS U2427 (.Y(n6559), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[12] ), 
	.B0(FE_OFN389_n4730), 
	.A1(FE_OFN1738_acc_fir_data_in_12_), 
	.A0(FE_OFN617_n4729));
   AO22XLTS U2413 (.Y(n6545), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[26] ), 
	.B0(FE_OFN386_n4730), 
	.A1(FE_OFN1659_acc_fir_data_in_26_), 
	.A0(FE_OFN611_n4729));
   AO22XLTS U2414 (.Y(n6546), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[25] ), 
	.B0(FE_OFN385_n4730), 
	.A1(FE_OFN1662_acc_fir_data_in_25_), 
	.A0(FE_OFN612_n4729));
   AO22XLTS U2424 (.Y(n6556), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[15] ), 
	.B0(FE_OFN389_n4730), 
	.A1(FE_OFN1720_acc_fir_data_in_15_), 
	.A0(FE_OFN617_n4729));
   AO22XLTS U2415 (.Y(n6547), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[24] ), 
	.B0(FE_OFN385_n4730), 
	.A1(FE_OFN1667_acc_fir_data_in_24_), 
	.A0(FE_OFN612_n4729));
   AO22XLTS U2412 (.Y(n6544), 
	.B1(\fifo_from_fir/fifo_cell6/sr_out[27] ), 
	.B0(FE_OFN386_n4730), 
	.A1(FE_OFN1652_acc_fir_data_in_27_), 
	.A0(FE_OFN611_n4729));
   AO22XLTS U1808 (.Y(n6042), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[0] ), 
	.B0(FE_OFN262_n4544), 
	.A1(FE_OFN1626_acc_fft_data_in_0_), 
	.A0(FE_OFN278_n4543));
   AO22XLTS U1797 (.Y(n6031), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[11] ), 
	.B0(FE_OFN261_n4544), 
	.A1(FE_OFN1563_acc_fft_data_in_11_), 
	.A0(FE_OFN272_n4543));
   AO22XLTS U1798 (.Y(n6032), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[10] ), 
	.B0(FE_OFN265_n4544), 
	.A1(FE_OFN1566_acc_fft_data_in_10_), 
	.A0(FE_OFN275_n4543));
   AO22XLTS U1795 (.Y(n6029), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[13] ), 
	.B0(FE_OFN261_n4544), 
	.A1(FE_OFN1548_acc_fft_data_in_13_), 
	.A0(FE_OFN272_n4543));
   AO22XLTS U1799 (.Y(n6033), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[9] ), 
	.B0(FE_OFN261_n4544), 
	.A1(FE_OFN1569_acc_fft_data_in_9_), 
	.A0(FE_OFN272_n4543));
   OAI21XLTS U845 (.Y(n3910), 
	.B0(n3912), 
	.A1(n3908), 
	.A0(n7276));
   AO22XLTS U1784 (.Y(n6018), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[24] ), 
	.B0(FE_OFN258_n4544), 
	.A1(FE_OFN1492_acc_fft_data_in_24_), 
	.A0(FE_OFN273_n4543));
   AO22XLTS U1807 (.Y(n6041), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[1] ), 
	.B0(FE_OFN259_n4544), 
	.A1(FE_OFN1620_acc_fft_data_in_1_), 
	.A0(FE_OFN276_n4543));
   AO22XLTS U1793 (.Y(n6027), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[15] ), 
	.B0(FE_OFN260_n4544), 
	.A1(FE_OFN1538_acc_fft_data_in_15_), 
	.A0(FE_OFN268_n4543));
   OAI21XLTS U989 (.Y(n4085), 
	.B0(n4087), 
	.A1(n4083), 
	.A0(n7385));
   AO22XLTS U1783 (.Y(n6017), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[25] ), 
	.B0(FE_OFN258_n4544), 
	.A1(FE_OFN1487_acc_fft_data_in_25_), 
	.A0(FE_OFN273_n4543));
   AO22XLTS U1782 (.Y(n6016), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[26] ), 
	.B0(FE_OFN262_n4544), 
	.A1(FE_OFN1482_acc_fft_data_in_26_), 
	.A0(FE_OFN278_n4543));
   AO22XLTS U1801 (.Y(n6035), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[7] ), 
	.B0(FE_OFN258_n4544), 
	.A1(FE_OFN1584_acc_fft_data_in_7_), 
	.A0(FE_OFN270_n4543));
   AO22XLTS U1802 (.Y(n6036), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[6] ), 
	.B0(FE_OFN256_n4544), 
	.A1(FE_OFN1589_acc_fft_data_in_6_), 
	.A0(FE_OFN269_n4543));
   AO22XLTS U1794 (.Y(n6028), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[14] ), 
	.B0(FE_OFN260_n4544), 
	.A1(FE_OFN1543_acc_fft_data_in_14_), 
	.A0(FE_OFN268_n4543));
   AO22XLTS U1806 (.Y(n6040), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[2] ), 
	.B0(FE_OFN259_n4544), 
	.A1(FE_OFN1614_acc_fft_data_in_2_), 
	.A0(FE_OFN276_n4543));
   AO22XLTS U1781 (.Y(n6015), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[27] ), 
	.B0(FE_OFN259_n4544), 
	.A1(FE_OFN1477_acc_fft_data_in_27_), 
	.A0(FE_OFN278_n4543));
   AO22XLTS U1800 (.Y(n6034), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[8] ), 
	.B0(FE_OFN261_n4544), 
	.A1(FE_OFN1575_acc_fft_data_in_8_), 
	.A0(FE_OFN272_n4543));
   AO22XLTS U1796 (.Y(n6030), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[12] ), 
	.B0(FE_OFN260_n4544), 
	.A1(FE_OFN1553_acc_fft_data_in_12_), 
	.A0(FE_OFN268_n4543));
   AO22XLTS U1805 (.Y(n6039), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[3] ), 
	.B0(FE_OFN262_n4544), 
	.A1(FE_OFN1607_acc_fft_data_in_3_), 
	.A0(FE_OFN278_n4543));
   OAI21XLTS U2406 (.Y(n4725), 
	.B0(FE_OFN593_n4723), 
	.A1(n4728), 
	.A0(n7569));
   AO22XLTS U1803 (.Y(n6037), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[5] ), 
	.B0(FE_OFN263_n4544), 
	.A1(FE_OFN1592_acc_fft_data_in_5_), 
	.A0(FE_OFN271_n4543));
   AO22XLTS U1804 (.Y(n6038), 
	.B1(\fifo_from_fft/fifo_cell6/sr_out[4] ), 
	.B0(FE_OFN256_n4544), 
	.A1(FE_OFN1600_acc_fft_data_in_4_), 
	.A0(FE_OFN269_n4543));
   NAND3XLTS U2670 (.Y(n4657), 
	.C(n4808), 
	.B(n4658), 
	.A(FE_OFN593_n4723));
   OAI21XLTS U1775 (.Y(n4539), 
	.B0(FE_OFN247_n4537), 
	.A1(n4542), 
	.A0(n7494));
   NAND3XLTS U1050 (.Y(n4045), 
	.C(n4151), 
	.B(n4046), 
	.A(n4087));
   OAI21XLTS U986 (.Y(n5537), 
	.B0(n4085), 
	.A1(n4084), 
	.A0(\fifo_to_fir/fifo_cell10/data_out/N35 ));
   NAND3XLTS U906 (.Y(n3870), 
	.C(n3976), 
	.B(n3871), 
	.A(n3912));
   OAI21XLTS U2405 (.Y(n6539), 
	.B0(n4725), 
	.A1(n4727), 
	.A0(\fifo_from_fir/fifo_cell7/data_out/N35 ));
   AOI21X1TS U844 (.Y(n5486), 
	.B0(FE_OFN842_n7619), 
	.A1(n3910), 
	.A0(\fifo_to_fft/fifo_cell10/controller/valid_read ));
   OAI21XLTS U842 (.Y(n5485), 
	.B0(n3910), 
	.A1(n3909), 
	.A0(\fifo_to_fft/fifo_cell10/data_out/N35 ));
   AOI21X1TS U988 (.Y(n5538), 
	.B0(FE_OFN800_n7619), 
	.A1(n4085), 
	.A0(\fifo_to_fir/fifo_cell10/controller/valid_read ));
   AOI21X1TS U2404 (.Y(n6538), 
	.B0(FE_OFN829_n7619), 
	.A1(n4725), 
	.A0(\fifo_from_fir/fifo_cell7/controller/valid_read ));
   AO22XLTS U2372 (.Y(n6507), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[30] ), 
	.B0(FE_OFN586_n4724), 
	.A1(FE_OFN1636_acc_fir_data_in_30_), 
	.A0(FE_OFN600_n4723));
   AO22XLTS U2371 (.Y(n6506), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[31] ), 
	.B0(FE_OFN588_n4724), 
	.A1(FE_OFN1628_acc_fir_data_in_31_), 
	.A0(FE_OFN599_n4723));
   OAI211XLTS U2671 (.Y(n4807), 
	.C0(n9467), 
	.B0(\fifo_from_fir/hang[6] ), 
	.A1(n4809), 
	.A0(n8875));
   AO22XLTS U2387 (.Y(n6522), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[15] ), 
	.B0(FE_OFN592_n4724), 
	.A1(FE_OFN1720_acc_fir_data_in_15_), 
	.A0(FE_OFN605_n4723));
   AO22XLTS U2373 (.Y(n6508), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[29] ), 
	.B0(FE_OFN588_n4724), 
	.A1(FE_OFN1640_acc_fir_data_in_29_), 
	.A0(FE_OFN599_n4723));
   AOI21X1TS U1773 (.Y(n6009), 
	.B0(FE_OFN825_n7619), 
	.A1(n4539), 
	.A0(\fifo_from_fft/fifo_cell7/controller/valid_read ));
   OAI211XLTS U907 (.Y(n3975), 
	.C0(n9479), 
	.B0(\fifo_to_fft/hang[9] ), 
	.A1(n3977), 
	.A0(n8809));
   AO22XLTS U2388 (.Y(n6523), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[14] ), 
	.B0(FE_OFN592_n4724), 
	.A1(FE_OFN1725_acc_fir_data_in_14_), 
	.A0(FE_OFN605_n4723));
   NAND3XLTS U2039 (.Y(n4471), 
	.C(n4622), 
	.B(n4472), 
	.A(FE_OFN250_n4537));
   AO22XLTS U2389 (.Y(n6524), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[13] ), 
	.B0(FE_OFN587_n4724), 
	.A1(FE_OFN1732_acc_fir_data_in_13_), 
	.A0(FE_OFN601_n4723));
   AO22XLTS U2390 (.Y(n6525), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[12] ), 
	.B0(FE_OFN592_n4724), 
	.A1(FE_OFN1738_acc_fir_data_in_12_), 
	.A0(FE_OFN605_n4723));
   OAI211XLTS U1051 (.Y(n4150), 
	.C0(n9475), 
	.B0(\fifo_to_fir/hang[9] ), 
	.A1(n4152), 
	.A0(n8788));
   AO22XLTS U2374 (.Y(n6509), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[28] ), 
	.B0(FE_OFN588_n4724), 
	.A1(FE_OFN1649_acc_fir_data_in_28_), 
	.A0(FE_OFN599_n4723));
   OAI21XLTS U1774 (.Y(n6010), 
	.B0(n4539), 
	.A1(n4541), 
	.A0(\fifo_from_fft/fifo_cell7/data_out/N35 ));
   AO22XLTS U1743 (.Y(n5980), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[28] ), 
	.B0(FE_OFN51_n4538), 
	.A1(FE_OFN1468_acc_fft_data_in_28_), 
	.A0(FE_OFN254_n4537));
   AO22XLTS U2401 (.Y(n6536), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[1] ), 
	.B0(n4724), 
	.A1(FE_OFN1807_acc_fir_data_in_1_), 
	.A0(n4723));
   AO22XLTS U1741 (.Y(n5978), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[30] ), 
	.B0(FE_OFN49_n4538), 
	.A1(FE_OFN1460_acc_fft_data_in_30_), 
	.A0(FE_OFN253_n4537));
   AO22XLTS U1740 (.Y(n5977), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[31] ), 
	.B0(FE_OFN49_n4538), 
	.A1(FE_OFN1455_acc_fft_data_in_31_), 
	.A0(FE_OFN253_n4537));
   OAI211XLTS U2040 (.Y(n4621), 
	.C0(n9471), 
	.B0(\fifo_from_fft/hang[6] ), 
	.A1(n4623), 
	.A0(n8842));
   AO22XLTS U2399 (.Y(n6534), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[3] ), 
	.B0(FE_OFN583_n4724), 
	.A1(FE_OFN1790_acc_fir_data_in_3_), 
	.A0(FE_OFN594_n4723));
   AO22XLTS U2384 (.Y(n6519), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[18] ), 
	.B0(FE_OFN587_n4724), 
	.A1(FE_OFN1702_acc_fir_data_in_18_), 
	.A0(FE_OFN601_n4723));
   AO22XLTS U2380 (.Y(n6515), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[22] ), 
	.B0(FE_OFN592_n4724), 
	.A1(FE_OFN1682_acc_fir_data_in_22_), 
	.A0(FE_OFN605_n4723));
   AO22XLTS U1756 (.Y(n5993), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[15] ), 
	.B0(FE_OFN48_n4538), 
	.A1(FE_OFN1541_acc_fft_data_in_15_), 
	.A0(FE_OFN246_n4537));
   AO22XLTS U2398 (.Y(n6533), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[4] ), 
	.B0(FE_OFN584_n4724), 
	.A1(FE_OFN1784_acc_fir_data_in_4_), 
	.A0(FE_OFN596_n4723));
   AO22XLTS U2375 (.Y(n6510), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[27] ), 
	.B0(FE_OFN590_n4724), 
	.A1(FE_OFN1652_acc_fir_data_in_27_), 
	.A0(FE_OFN600_n4723));
   AO22XLTS U2400 (.Y(n6535), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[2] ), 
	.B0(FE_OFN583_n4724), 
	.A1(FE_OFN1801_acc_fir_data_in_2_), 
	.A0(FE_OFN596_n4723));
   AO22XLTS U2385 (.Y(n6520), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[17] ), 
	.B0(FE_OFN585_n4724), 
	.A1(FE_OFN1707_acc_fir_data_in_17_), 
	.A0(FE_OFN598_n4723));
   AO22XLTS U2386 (.Y(n6521), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[16] ), 
	.B0(FE_OFN585_n4724), 
	.A1(FE_OFN1713_acc_fir_data_in_16_), 
	.A0(FE_OFN601_n4723));
   AO22XLTS U2397 (.Y(n6532), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[5] ), 
	.B0(FE_OFN584_n4724), 
	.A1(FE_OFN1778_acc_fir_data_in_5_), 
	.A0(FE_OFN597_n4723));
   AO22XLTS U2378 (.Y(n6513), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[24] ), 
	.B0(FE_OFN590_n4724), 
	.A1(FE_OFN1668_acc_fir_data_in_24_), 
	.A0(FE_OFN602_n4723));
   AO22XLTS U1759 (.Y(n5996), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[12] ), 
	.B0(FE_OFN46_n4538), 
	.A1(FE_OFN1558_acc_fft_data_in_12_), 
	.A0(FE_OFN244_n4537));
   AO22XLTS U2376 (.Y(n6511), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[26] ), 
	.B0(FE_OFN590_n4724), 
	.A1(FE_OFN1660_acc_fir_data_in_26_), 
	.A0(FE_OFN600_n4723));
   AO22XLTS U2379 (.Y(n6514), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[23] ), 
	.B0(FE_OFN585_n4724), 
	.A1(FE_OFN1675_acc_fir_data_in_23_), 
	.A0(FE_OFN598_n4723));
   AO22XLTS U2402 (.Y(n6537), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[0] ), 
	.B0(FE_OFN583_n4724), 
	.A1(FE_OFN1813_acc_fir_data_in_0_), 
	.A0(FE_OFN594_n4723));
   AO22XLTS U2396 (.Y(n6531), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[6] ), 
	.B0(FE_OFN586_n4724), 
	.A1(FE_OFN1771_acc_fir_data_in_6_), 
	.A0(FE_OFN597_n4723));
   AO22XLTS U2383 (.Y(n6518), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[19] ), 
	.B0(FE_OFN582_n4724), 
	.A1(FE_OFN1700_acc_fir_data_in_19_), 
	.A0(FE_OFN595_n4723));
   AO22XLTS U2394 (.Y(n6529), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[8] ), 
	.B0(FE_OFN589_n4724), 
	.A1(FE_OFN1756_acc_fir_data_in_8_), 
	.A0(FE_OFN604_n4723));
   AO22XLTS U2381 (.Y(n6516), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[21] ), 
	.B0(FE_OFN582_n4724), 
	.A1(FE_OFN1687_acc_fir_data_in_21_), 
	.A0(FE_OFN598_n4723));
   AO22XLTS U2393 (.Y(n6528), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[9] ), 
	.B0(FE_OFN589_n4724), 
	.A1(FE_OFN1752_acc_fir_data_in_9_), 
	.A0(FE_OFN604_n4723));
   AO22XLTS U2395 (.Y(n6530), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[7] ), 
	.B0(FE_OFN584_n4724), 
	.A1(FE_OFN1766_acc_fir_data_in_7_), 
	.A0(FE_OFN596_n4723));
   AO22XLTS U2377 (.Y(n6512), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[25] ), 
	.B0(FE_OFN590_n4724), 
	.A1(FE_OFN1663_acc_fir_data_in_25_), 
	.A0(FE_OFN602_n4723));
   AO22XLTS U2392 (.Y(n6527), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[10] ), 
	.B0(FE_OFN591_n4724), 
	.A1(FE_OFN1747_acc_fir_data_in_10_), 
	.A0(FE_OFN603_n4723));
   AO22XLTS U2382 (.Y(n6517), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[20] ), 
	.B0(FE_OFN582_n4724), 
	.A1(FE_OFN1693_acc_fir_data_in_20_), 
	.A0(FE_OFN595_n4723));
   AO22XLTS U2391 (.Y(n6526), 
	.B1(\fifo_from_fir/fifo_cell7/sr_out[11] ), 
	.B0(FE_OFN589_n4724), 
	.A1(FE_OFN1745_acc_fir_data_in_11_), 
	.A0(FE_OFN604_n4723));
   AO22XLTS U1758 (.Y(n5995), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[13] ), 
	.B0(FE_OFN48_n4538), 
	.A1(FE_OFN1551_acc_fft_data_in_13_), 
	.A0(FE_OFN246_n4537));
   AO22XLTS U1742 (.Y(n5979), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[29] ), 
	.B0(FE_OFN49_n4538), 
	.A1(FE_OFN1464_acc_fft_data_in_29_), 
	.A0(FE_OFN253_n4537));
   AO22XLTS U1757 (.Y(n5994), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[14] ), 
	.B0(FE_OFN48_n4538), 
	.A1(FE_OFN1547_acc_fft_data_in_14_), 
	.A0(FE_OFN246_n4537));
   AO22XLTS U1746 (.Y(n5983), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[25] ), 
	.B0(FE_OFN44_n4538), 
	.A1(FE_OFN1485_acc_fft_data_in_25_), 
	.A0(FE_OFN248_n4537));
   AO22XLTS U1766 (.Y(n6003), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[5] ), 
	.B0(FE_OFN45_n4538), 
	.A1(FE_OFN1594_acc_fft_data_in_5_), 
	.A0(FE_OFN251_n4537));
   AO22XLTS U1763 (.Y(n6000), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[8] ), 
	.B0(FE_OFN52_n4538), 
	.A1(FE_OFN1577_acc_fft_data_in_8_), 
	.A0(FE_OFN255_n4537));
   NAND3XLTS U904 (.Y(n3872), 
	.C(n3973), 
	.B(n3873), 
	.A(n3907));
   AO22XLTS U1765 (.Y(n6002), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[6] ), 
	.B0(FE_OFN50_n4538), 
	.A1(FE_OFN1587_acc_fft_data_in_6_), 
	.A0(FE_OFN249_n4537));
   AO22XLTS U1744 (.Y(n5981), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[27] ), 
	.B0(FE_OFN45_n4538), 
	.A1(FE_OFN1476_acc_fft_data_in_27_), 
	.A0(FE_OFN251_n4537));
   AO22XLTS U1769 (.Y(n6006), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[2] ), 
	.B0(FE_OFN44_n4538), 
	.A1(FE_OFN1612_acc_fft_data_in_2_), 
	.A0(FE_OFN248_n4537));
   AO22XLTS U1761 (.Y(n5998), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[10] ), 
	.B0(FE_OFN52_n4538), 
	.A1(FE_OFN1565_acc_fft_data_in_10_), 
	.A0(FE_OFN255_n4537));
   AO22XLTS U1760 (.Y(n5997), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[11] ), 
	.B0(FE_OFN52_n4538), 
	.A1(FE_OFN1561_acc_fft_data_in_11_), 
	.A0(FE_OFN255_n4537));
   AO22XLTS U1748 (.Y(n5985), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[23] ), 
	.B0(FE_OFN50_n4538), 
	.A1(FE_OFN1497_acc_fft_data_in_23_), 
	.A0(FE_OFN249_n4537));
   AO22XLTS U1768 (.Y(n6005), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[3] ), 
	.B0(FE_OFN47_n4538), 
	.A1(FE_OFN1606_acc_fft_data_in_3_), 
	.A0(FE_OFN252_n4537));
   AO22XLTS U1762 (.Y(n5999), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[9] ), 
	.B0(FE_OFN52_n4538), 
	.A1(FE_OFN1573_acc_fft_data_in_9_), 
	.A0(FE_OFN255_n4537));
   AO22XLTS U1750 (.Y(n5987), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[21] ), 
	.B0(FE_OFN51_n4538), 
	.A1(FE_OFN1507_acc_fft_data_in_21_), 
	.A0(FE_OFN254_n4537));
   AO22XLTS U1749 (.Y(n5986), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[22] ), 
	.B0(FE_OFN51_n4538), 
	.A1(FE_OFN1500_acc_fft_data_in_22_), 
	.A0(FE_OFN254_n4537));
   AO22XLTS U1770 (.Y(n6007), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[1] ), 
	.B0(FE_OFN45_n4538), 
	.A1(FE_OFN1618_acc_fft_data_in_1_), 
	.A0(FE_OFN251_n4537));
   AO22XLTS U1745 (.Y(n5982), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[26] ), 
	.B0(FE_OFN47_n4538), 
	.A1(FE_OFN1480_acc_fft_data_in_26_), 
	.A0(FE_OFN252_n4537));
   AO22XLTS U1747 (.Y(n5984), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[24] ), 
	.B0(FE_OFN44_n4538), 
	.A1(FE_OFN1491_acc_fft_data_in_24_), 
	.A0(FE_OFN250_n4537));
   NAND3XLTS U1048 (.Y(n4047), 
	.C(n4148), 
	.B(n4048), 
	.A(n4082));
   AO22XLTS U1751 (.Y(n5988), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[20] ), 
	.B0(FE_OFN50_n4538), 
	.A1(FE_OFN1512_acc_fft_data_in_20_), 
	.A0(FE_OFN249_n4537));
   AO22XLTS U1752 (.Y(n5989), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[19] ), 
	.B0(FE_OFN43_n4538), 
	.A1(FE_OFN1519_acc_fft_data_in_19_), 
	.A0(n4537));
   AO22XLTS U1753 (.Y(n5990), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[18] ), 
	.B0(FE_OFN50_n4538), 
	.A1(FE_OFN1523_acc_fft_data_in_18_), 
	.A0(FE_OFN249_n4537));
   AO22XLTS U1767 (.Y(n6004), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[4] ), 
	.B0(FE_OFN43_n4538), 
	.A1(FE_OFN1599_acc_fft_data_in_4_), 
	.A0(FE_OFN245_n4537));
   AO22XLTS U1754 (.Y(n5991), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[17] ), 
	.B0(FE_OFN46_n4538), 
	.A1(FE_OFN1531_acc_fft_data_in_17_), 
	.A0(FE_OFN244_n4537));
   AO22XLTS U1764 (.Y(n6001), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[7] ), 
	.B0(n4538), 
	.A1(FE_OFN1584_acc_fft_data_in_7_), 
	.A0(FE_OFN245_n4537));
   AO22XLTS U1755 (.Y(n5992), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[16] ), 
	.B0(FE_OFN46_n4538), 
	.A1(FE_OFN1536_acc_fft_data_in_16_), 
	.A0(n4537));
   AO22XLTS U1771 (.Y(n6008), 
	.B1(\fifo_from_fft/fifo_cell7/sr_out[0] ), 
	.B0(FE_OFN47_n4538), 
	.A1(FE_OFN1624_acc_fft_data_in_0_), 
	.A0(FE_OFN252_n4537));
   OAI211XLTS U1049 (.Y(n4147), 
	.C0(n9475), 
	.B0(\fifo_to_fir/hang[10] ), 
	.A1(n4149), 
	.A0(n8788));
   OAI211XLTS U905 (.Y(n3972), 
	.C0(n9479), 
	.B0(\fifo_to_fft/hang[10] ), 
	.A1(n3974), 
	.A0(n8809));
   OAI21XLTS U2369 (.Y(n4719), 
	.B0(n4717), 
	.A1(n4722), 
	.A0(n7564));
   OAI21XLTS U1738 (.Y(n4533), 
	.B0(FE_OFN233_n4531), 
	.A1(n4536), 
	.A0(n7490));
   OAI21XLTS U2368 (.Y(n6505), 
	.B0(n4719), 
	.A1(n4721), 
	.A0(\fifo_from_fir/fifo_cell8/data_out/N35 ));
   NAND3XLTS U2668 (.Y(n4659), 
	.C(n4805), 
	.B(n4660), 
	.A(n4717));
   AO22XLTS U2343 (.Y(n6481), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[22] ), 
	.B0(FE_OFN400_n4718), 
	.A1(FE_OFN1680_acc_fir_data_in_22_), 
	.A0(FE_OFN577_n4717));
   AOI21X1TS U2367 (.Y(n6504), 
	.B0(FE_OFN817_n7619), 
	.A1(n4719), 
	.A0(\fifo_from_fir/fifo_cell8/controller/valid_read ));
   AO22XLTS U2344 (.Y(n6482), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[21] ), 
	.B0(FE_OFN396_n4718), 
	.A1(FE_OFN1689_acc_fir_data_in_21_), 
	.A0(FE_OFN573_n4717));
   NAND3XLTS U2037 (.Y(n4473), 
	.C(n4619), 
	.B(n4474), 
	.A(n4531));
   AO22XLTS U1713 (.Y(n5953), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[21] ), 
	.B0(FE_OFN57_n4532), 
	.A1(FE_OFN1506_acc_fft_data_in_21_), 
	.A0(FE_OFN239_n4531));
   AO22XLTS U1712 (.Y(n5952), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[22] ), 
	.B0(FE_OFN57_n4532), 
	.A1(FE_OFN1504_acc_fft_data_in_22_), 
	.A0(FE_OFN239_n4531));
   OAI21XLTS U1737 (.Y(n5976), 
	.B0(n4533), 
	.A1(n4535), 
	.A0(\fifo_from_fft/fifo_cell8/data_out/N35 ));
   AOI21X1TS U1736 (.Y(n5975), 
	.B0(FE_OFN827_n7619), 
	.A1(n4533), 
	.A0(\fifo_from_fft/fifo_cell8/controller/valid_read ));
   AO22XLTS U2334 (.Y(n6472), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[31] ), 
	.B0(FE_OFN399_n4718), 
	.A1(FE_OFN1629_acc_fir_data_in_31_), 
	.A0(FE_OFN581_n4717));
   AO22XLTS U2336 (.Y(n6474), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[29] ), 
	.B0(FE_OFN399_n4718), 
	.A1(FE_OFN1641_acc_fir_data_in_29_), 
	.A0(FE_OFN581_n4717));
   OAI211XLTS U2669 (.Y(n4804), 
	.C0(n9467), 
	.B0(\fifo_from_fir/hang[7] ), 
	.A1(n4806), 
	.A0(n8875));
   AO22XLTS U2342 (.Y(n6480), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[23] ), 
	.B0(FE_OFN396_n4718), 
	.A1(FE_OFN1676_acc_fir_data_in_23_), 
	.A0(FE_OFN573_n4717));
   AO22XLTS U2335 (.Y(n6473), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[30] ), 
	.B0(FE_OFN399_n4718), 
	.A1(FE_OFN1634_acc_fir_data_in_30_), 
	.A0(FE_OFN581_n4717));
   AO22XLTS U2345 (.Y(n6483), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[20] ), 
	.B0(n4718), 
	.A1(FE_OFN1692_acc_fir_data_in_20_), 
	.A0(FE_OFN571_n4717));
   AO22XLTS U2346 (.Y(n6484), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[19] ), 
	.B0(FE_OFN393_n4718), 
	.A1(FE_OFN1695_acc_fir_data_in_19_), 
	.A0(FE_OFN574_n4717));
   NAND3XLTS U902 (.Y(n3874), 
	.C(n3970), 
	.B(n3875), 
	.A(n7265));
   AO22XLTS U2349 (.Y(n6487), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[16] ), 
	.B0(FE_OFN394_n4718), 
	.A1(FE_OFN1716_acc_fir_data_in_16_), 
	.A0(FE_OFN576_n4717));
   AO22XLTS U2347 (.Y(n6485), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[18] ), 
	.B0(FE_OFN394_n4718), 
	.A1(FE_OFN1702_acc_fir_data_in_18_), 
	.A0(FE_OFN576_n4717));
   AO22XLTS U1703 (.Y(n5943), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[31] ), 
	.B0(FE_OFN55_n4532), 
	.A1(FE_OFN1456_acc_fft_data_in_31_), 
	.A0(FE_OFN240_n4531));
   AO22XLTS U1711 (.Y(n5951), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[23] ), 
	.B0(FE_OFN53_n4532), 
	.A1(FE_OFN1496_acc_fft_data_in_23_), 
	.A0(FE_OFN236_n4531));
   AO22XLTS U2348 (.Y(n6486), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[17] ), 
	.B0(FE_OFN393_n4718), 
	.A1(FE_OFN1707_acc_fir_data_in_17_), 
	.A0(FE_OFN576_n4717));
   AO22XLTS U1704 (.Y(n5944), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[30] ), 
	.B0(FE_OFN58_n4532), 
	.A1(FE_OFN1459_acc_fft_data_in_30_), 
	.A0(FE_OFN240_n4531));
   AO22XLTS U1714 (.Y(n5954), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[20] ), 
	.B0(FE_OFN54_n4532), 
	.A1(FE_OFN1512_acc_fft_data_in_20_), 
	.A0(FE_OFN238_n4531));
   AO22XLTS U1705 (.Y(n5945), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[29] ), 
	.B0(FE_OFN58_n4532), 
	.A1(FE_OFN1465_acc_fft_data_in_29_), 
	.A0(FE_OFN240_n4531));
   NAND3XLTS U1046 (.Y(n4049), 
	.C(n4145), 
	.B(n4050), 
	.A(n7374));
   OAI211XLTS U2038 (.Y(n4618), 
	.C0(n9471), 
	.B0(\fifo_from_fft/hang[7] ), 
	.A1(n4620), 
	.A0(n8842));
   AO22XLTS U2337 (.Y(n6475), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[28] ), 
	.B0(FE_OFN399_n4718), 
	.A1(FE_OFN1647_acc_fir_data_in_28_), 
	.A0(FE_OFN581_n4717));
   AO22XLTS U1716 (.Y(n5956), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[18] ), 
	.B0(FE_OFN54_n4532), 
	.A1(FE_OFN1523_acc_fft_data_in_18_), 
	.A0(FE_OFN238_n4531));
   AO22XLTS U2351 (.Y(n6489), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[14] ), 
	.B0(FE_OFN400_n4718), 
	.A1(FE_OFN1728_acc_fir_data_in_14_), 
	.A0(FE_OFN577_n4717));
   AO22XLTS U2365 (.Y(n6503), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[0] ), 
	.B0(FE_OFN393_n4718), 
	.A1(FE_OFN1817_acc_fir_data_in_0_), 
	.A0(FE_OFN574_n4717));
   AO22XLTS U2340 (.Y(n6478), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[25] ), 
	.B0(FE_OFN398_n4718), 
	.A1(FE_OFN1663_acc_fir_data_in_25_), 
	.A0(FE_OFN580_n4717));
   AO22XLTS U2353 (.Y(n6491), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[12] ), 
	.B0(FE_OFN400_n4718), 
	.A1(FE_OFN1737_acc_fir_data_in_12_), 
	.A0(FE_OFN577_n4717));
   AO22XLTS U2350 (.Y(n6488), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[15] ), 
	.B0(FE_OFN396_n4718), 
	.A1(FE_OFN1721_acc_fir_data_in_15_), 
	.A0(FE_OFN573_n4717));
   AO22XLTS U2355 (.Y(n6493), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[10] ), 
	.B0(FE_OFN400_n4718), 
	.A1(FE_OFN1748_acc_fir_data_in_10_), 
	.A0(FE_OFN577_n4717));
   AO22XLTS U1706 (.Y(n5946), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[28] ), 
	.B0(FE_OFN55_n4532), 
	.A1(FE_OFN1820_acc_fft_data_in_28_), 
	.A0(FE_OFN240_n4531));
   AO22XLTS U2364 (.Y(n6502), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[1] ), 
	.B0(FE_OFN391_n4718), 
	.A1(FE_OFN1807_acc_fir_data_in_1_), 
	.A0(FE_OFN570_n4717));
   AO22XLTS U2352 (.Y(n6490), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[13] ), 
	.B0(FE_OFN397_n4718), 
	.A1(FE_OFN1731_acc_fir_data_in_13_), 
	.A0(FE_OFN579_n4717));
   AO22XLTS U2363 (.Y(n6501), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[2] ), 
	.B0(FE_OFN392_n4718), 
	.A1(FE_OFN1796_acc_fir_data_in_2_), 
	.A0(FE_OFN572_n4717));
   AO22XLTS U2357 (.Y(n6495), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[8] ), 
	.B0(FE_OFN397_n4718), 
	.A1(FE_OFN1757_acc_fir_data_in_8_), 
	.A0(FE_OFN579_n4717));
   AO22XLTS U2354 (.Y(n6492), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[11] ), 
	.B0(FE_OFN397_n4718), 
	.A1(FE_OFN1741_acc_fir_data_in_11_), 
	.A0(FE_OFN579_n4717));
   AO22XLTS U2362 (.Y(n6500), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[3] ), 
	.B0(FE_OFN390_n4718), 
	.A1(FE_OFN1791_acc_fir_data_in_3_), 
	.A0(FE_OFN570_n4717));
   AO22XLTS U1715 (.Y(n5955), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[19] ), 
	.B0(FE_OFN59_n4532), 
	.A1(FE_OFN1519_acc_fft_data_in_19_), 
	.A0(FE_OFN243_n4531));
   AO22XLTS U1718 (.Y(n5958), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[16] ), 
	.B0(FE_OFN59_n4532), 
	.A1(FE_OFN1537_acc_fft_data_in_16_), 
	.A0(FE_OFN243_n4531));
   AO22XLTS U2339 (.Y(n6477), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[26] ), 
	.B0(FE_OFN398_n4718), 
	.A1(FE_OFN1659_acc_fir_data_in_26_), 
	.A0(FE_OFN578_n4717));
   OAI211XLTS U1047 (.Y(n4144), 
	.C0(n9476), 
	.B0(\fifo_to_fir/hang[11] ), 
	.A1(n4146), 
	.A0(n8788));
   AO22XLTS U2338 (.Y(n6476), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[27] ), 
	.B0(FE_OFN395_n4718), 
	.A1(FE_OFN1652_acc_fir_data_in_27_), 
	.A0(FE_OFN578_n4717));
   AO22XLTS U2356 (.Y(n6494), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[9] ), 
	.B0(FE_OFN397_n4718), 
	.A1(FE_OFN1751_acc_fir_data_in_9_), 
	.A0(FE_OFN579_n4717));
   AO22XLTS U2361 (.Y(n6499), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[4] ), 
	.B0(FE_OFN391_n4718), 
	.A1(FE_OFN1788_acc_fir_data_in_4_), 
	.A0(FE_OFN575_n4717));
   AO22XLTS U1717 (.Y(n5957), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[17] ), 
	.B0(FE_OFN59_n4532), 
	.A1(FE_OFN1532_acc_fft_data_in_17_), 
	.A0(FE_OFN243_n4531));
   AO22XLTS U2341 (.Y(n6479), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[24] ), 
	.B0(FE_OFN398_n4718), 
	.A1(FE_OFN1667_acc_fir_data_in_24_), 
	.A0(FE_OFN580_n4717));
   OAI211XLTS U903 (.Y(n3969), 
	.C0(n9479), 
	.B0(\fifo_to_fft/hang[11] ), 
	.A1(n3971), 
	.A0(n8809));
   AO22XLTS U2360 (.Y(n6498), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[5] ), 
	.B0(FE_OFN395_n4718), 
	.A1(FE_OFN1782_acc_fir_data_in_5_), 
	.A0(FE_OFN575_n4717));
   AO22XLTS U2358 (.Y(n6496), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[7] ), 
	.B0(FE_OFN392_n4718), 
	.A1(FE_OFN1763_acc_fir_data_in_7_), 
	.A0(FE_OFN572_n4717));
   AO22XLTS U2359 (.Y(n6497), 
	.B1(\fifo_from_fir/fifo_cell8/sr_out[6] ), 
	.B0(FE_OFN392_n4718), 
	.A1(FE_OFN1769_acc_fir_data_in_6_), 
	.A0(FE_OFN575_n4717));
   AO22XLTS U1734 (.Y(n5974), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[0] ), 
	.B0(FE_OFN58_n4532), 
	.A1(FE_OFN1626_acc_fft_data_in_0_), 
	.A0(FE_OFN237_n4531));
   AO22XLTS U1726 (.Y(n5966), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[8] ), 
	.B0(FE_OFN60_n4532), 
	.A1(FE_OFN1577_acc_fft_data_in_8_), 
	.A0(FE_OFN241_n4531));
   AO22XLTS U1728 (.Y(n5968), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[6] ), 
	.B0(FE_OFN53_n4532), 
	.A1(FE_OFN1588_acc_fft_data_in_6_), 
	.A0(FE_OFN235_n4531));
   AO22XLTS U1724 (.Y(n5964), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[10] ), 
	.B0(FE_OFN60_n4532), 
	.A1(FE_OFN1566_acc_fft_data_in_10_), 
	.A0(FE_OFN241_n4531));
   AO22XLTS U1730 (.Y(n5970), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[4] ), 
	.B0(n4532), 
	.A1(FE_OFN1602_acc_fft_data_in_4_), 
	.A0(FE_OFN235_n4531));
   AO22XLTS U1729 (.Y(n5969), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[5] ), 
	.B0(n4532), 
	.A1(FE_OFN1594_acc_fft_data_in_5_), 
	.A0(FE_OFN236_n4531));
   AO22XLTS U1731 (.Y(n5971), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[3] ), 
	.B0(FE_OFN61_n4532), 
	.A1(FE_OFN1607_acc_fft_data_in_3_), 
	.A0(FE_OFN237_n4531));
   AO22XLTS U1719 (.Y(n5959), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[15] ), 
	.B0(FE_OFN56_n4532), 
	.A1(FE_OFN1540_acc_fft_data_in_15_), 
	.A0(FE_OFN242_n4531));
   AO22XLTS U1722 (.Y(n5962), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[12] ), 
	.B0(FE_OFN59_n4532), 
	.A1(FE_OFN1558_acc_fft_data_in_12_), 
	.A0(FE_OFN243_n4531));
   AO22XLTS U1732 (.Y(n5972), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[2] ), 
	.B0(FE_OFN62_n4532), 
	.A1(FE_OFN1614_acc_fft_data_in_2_), 
	.A0(FE_OFN234_n4531));
   AO22XLTS U1727 (.Y(n5967), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[7] ), 
	.B0(n4532), 
	.A1(FE_OFN1582_acc_fft_data_in_7_), 
	.A0(FE_OFN235_n4531));
   AO22XLTS U1723 (.Y(n5963), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[11] ), 
	.B0(FE_OFN60_n4532), 
	.A1(FE_OFN1562_acc_fft_data_in_11_), 
	.A0(FE_OFN241_n4531));
   AO22XLTS U1721 (.Y(n5961), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[13] ), 
	.B0(FE_OFN56_n4532), 
	.A1(FE_OFN1552_acc_fft_data_in_13_), 
	.A0(FE_OFN242_n4531));
   AO22XLTS U1720 (.Y(n5960), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[14] ), 
	.B0(FE_OFN56_n4532), 
	.A1(FE_OFN1547_acc_fft_data_in_14_), 
	.A0(FE_OFN242_n4531));
   AO22XLTS U1725 (.Y(n5965), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[9] ), 
	.B0(FE_OFN60_n4532), 
	.A1(FE_OFN1572_acc_fft_data_in_9_), 
	.A0(FE_OFN241_n4531));
   AO22XLTS U1733 (.Y(n5973), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[1] ), 
	.B0(FE_OFN62_n4532), 
	.A1(FE_OFN1620_acc_fft_data_in_1_), 
	.A0(FE_OFN234_n4531));
   AO22XLTS U1710 (.Y(n5950), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[24] ), 
	.B0(FE_OFN62_n4532), 
	.A1(FE_OFN1491_acc_fft_data_in_24_), 
	.A0(FE_OFN232_n4531));
   AO22XLTS U1709 (.Y(n5949), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[25] ), 
	.B0(FE_OFN62_n4532), 
	.A1(FE_OFN1487_acc_fft_data_in_25_), 
	.A0(FE_OFN234_n4531));
   AO22XLTS U1707 (.Y(n5947), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[27] ), 
	.B0(FE_OFN61_n4532), 
	.A1(FE_OFN1477_acc_fft_data_in_27_), 
	.A0(FE_OFN237_n4531));
   AO22XLTS U1708 (.Y(n5948), 
	.B1(\fifo_from_fft/fifo_cell8/sr_out[26] ), 
	.B0(FE_OFN61_n4532), 
	.A1(FE_OFN1482_acc_fft_data_in_26_), 
	.A0(FE_OFN237_n4531));
   OAI21XLTS U2332 (.Y(n4713), 
	.B0(n4711), 
	.A1(n4716), 
	.A0(n7559));
   NAND3XLTS U2666 (.Y(n4661), 
	.C(n4802), 
	.B(n4662), 
	.A(n4711));
   OAI21XLTS U2331 (.Y(n6471), 
	.B0(n4713), 
	.A1(n4715), 
	.A0(\fifo_from_fir/fifo_cell9/data_out/N35 ));
   OAI21X1TS U1701 (.Y(n4527), 
	.B0(n4525), 
	.A1(n4530), 
	.A0(n7485));
   AO22XLTS U2322 (.Y(n6463), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[6] ), 
	.B0(FE_OFN427_n4712), 
	.A1(FE_OFN1773_acc_fir_data_in_6_), 
	.A0(FE_OFN561_n4711));
   AOI21X1TS U2330 (.Y(n6470), 
	.B0(FE_OFN817_n7619), 
	.A1(n4713), 
	.A0(\fifo_from_fir/fifo_cell9/controller/valid_read ));
   AO22XLTS U2297 (.Y(n6438), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[31] ), 
	.B0(FE_OFN430_n4712), 
	.A1(FE_OFN1628_acc_fir_data_in_31_), 
	.A0(FE_OFN567_n4711));
   OAI211XLTS U2667 (.Y(n4801), 
	.C0(n9467), 
	.B0(\fifo_from_fir/hang[8] ), 
	.A1(n4803), 
	.A0(n8875));
   AO22XLTS U2327 (.Y(n6468), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[1] ), 
	.B0(n4712), 
	.A1(FE_OFN1806_acc_fir_data_in_1_), 
	.A0(FE_OFN560_n4711));
   AO22XLTS U2326 (.Y(n6467), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[2] ), 
	.B0(FE_OFN425_n4712), 
	.A1(FE_OFN1796_acc_fir_data_in_2_), 
	.A0(FE_OFN561_n4711));
   AO22XLTS U2299 (.Y(n6440), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[29] ), 
	.B0(FE_OFN430_n4712), 
	.A1(FE_OFN1642_acc_fir_data_in_29_), 
	.A0(FE_OFN567_n4711));
   NAND3XLTS U2035 (.Y(n4475), 
	.C(n4616), 
	.B(n4476), 
	.A(FE_OFN221_n4525));
   AO22XLTS U2324 (.Y(n6465), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[4] ), 
	.B0(FE_OFN423_n4712), 
	.A1(FE_OFN1788_acc_fir_data_in_4_), 
	.A0(FE_OFN558_n4711));
   NAND3XLTS U900 (.Y(n3876), 
	.C(n3967), 
	.B(n3877), 
	.A(n7255));
   AO22XLTS U2323 (.Y(n6464), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[5] ), 
	.B0(FE_OFN427_n4712), 
	.A1(FE_OFN1782_acc_fir_data_in_5_), 
	.A0(FE_OFN564_n4711));
   OAI21XLTS U1700 (.Y(n5942), 
	.B0(n4527), 
	.A1(n4529), 
	.A0(\fifo_from_fft/fifo_cell9/data_out/N35 ));
   AO22XLTS U2328 (.Y(n6469), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[0] ), 
	.B0(FE_OFN423_n4712), 
	.A1(FE_OFN1817_acc_fir_data_in_0_), 
	.A0(FE_OFN562_n4711));
   AO22XLTS U2321 (.Y(n6462), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[7] ), 
	.B0(FE_OFN425_n4712), 
	.A1(FE_OFN1767_acc_fir_data_in_7_), 
	.A0(FE_OFN561_n4711));
   NAND3XLTS U1044 (.Y(n4051), 
	.C(n4142), 
	.B(n4052), 
	.A(n7365));
   AO22XLTS U2298 (.Y(n6439), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[30] ), 
	.B0(FE_OFN430_n4712), 
	.A1(FE_OFN1633_acc_fir_data_in_30_), 
	.A0(FE_OFN567_n4711));
   AO22XLTS U2325 (.Y(n6466), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[3] ), 
	.B0(FE_OFN423_n4712), 
	.A1(FE_OFN1791_acc_fir_data_in_3_), 
	.A0(FE_OFN559_n4711));
   AOI21X1TS U1699 (.Y(n5941), 
	.B0(FE_OFN830_n7619), 
	.A1(n4527), 
	.A0(\fifo_from_fft/fifo_cell9/controller/valid_read ));
   AO22XLTS U1675 (.Y(n5918), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[22] ), 
	.B0(FE_OFN91_n4526), 
	.A1(FE_OFN1500_acc_fft_data_in_22_), 
	.A0(FE_OFN227_n4525));
   AO22XLTS U1677 (.Y(n5920), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[20] ), 
	.B0(FE_OFN93_n4526), 
	.A1(FE_OFN1510_acc_fft_data_in_20_), 
	.A0(FE_OFN230_n4525));
   AO22XLTS U1676 (.Y(n5919), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[21] ), 
	.B0(FE_OFN91_n4526), 
	.A1(FE_OFN1505_acc_fft_data_in_21_), 
	.A0(FE_OFN227_n4525));
   AO22XLTS U1674 (.Y(n5917), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[23] ), 
	.B0(FE_OFN87_n4526), 
	.A1(FE_OFN1497_acc_fft_data_in_23_), 
	.A0(FE_OFN225_n4525));
   OAI211XLTS U2036 (.Y(n4615), 
	.C0(n9471), 
	.B0(\fifo_from_fft/hang[8] ), 
	.A1(n4617), 
	.A0(n8842));
   OAI211XLTS U901 (.Y(n3966), 
	.C0(n9478), 
	.B0(\fifo_to_fft/hang[12] ), 
	.A1(n3968), 
	.A0(n8809));
   AO22XLTS U2300 (.Y(n6441), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[28] ), 
	.B0(FE_OFN430_n4712), 
	.A1(FE_OFN1647_acc_fir_data_in_28_), 
	.A0(FE_OFN567_n4711));
   OAI211XLTS U1045 (.Y(n4141), 
	.C0(n9474), 
	.B0(\fifo_to_fir/hang[12] ), 
	.A1(n4143), 
	.A0(n8788));
   AO22XLTS U1669 (.Y(n5912), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[28] ), 
	.B0(FE_OFN87_n4526), 
	.A1(FE_OFN1470_acc_fft_data_in_28_), 
	.A0(FE_OFN228_n4525));
   AO22XLTS U1668 (.Y(n5911), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[29] ), 
	.B0(FE_OFN90_n4526), 
	.A1(FE_OFN1463_acc_fft_data_in_29_), 
	.A0(FE_OFN228_n4525));
   AO22XLTS U1667 (.Y(n5910), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[30] ), 
	.B0(FE_OFN90_n4526), 
	.A1(FE_OFN1458_acc_fft_data_in_30_), 
	.A0(FE_OFN228_n4525));
   AO22XLTS U1666 (.Y(n5909), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[31] ), 
	.B0(FE_OFN90_n4526), 
	.A1(FE_OFN1457_acc_fft_data_in_31_), 
	.A0(FE_OFN228_n4525));
   AO22XLTS U2311 (.Y(n6452), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[17] ), 
	.B0(FE_OFN426_n4712), 
	.A1(FE_OFN1709_acc_fir_data_in_17_), 
	.A0(FE_OFN562_n4711));
   AO22XLTS U2310 (.Y(n6451), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[18] ), 
	.B0(FE_OFN426_n4712), 
	.A1(FE_OFN1703_acc_fir_data_in_18_), 
	.A0(FE_OFN563_n4711));
   AO22XLTS U1687 (.Y(n5930), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[10] ), 
	.B0(FE_OFN91_n4526), 
	.A1(FE_OFN1564_acc_fft_data_in_10_), 
	.A0(FE_OFN229_n4525));
   AO22XLTS U1678 (.Y(n5921), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[19] ), 
	.B0(FE_OFN85_n4526), 
	.A1(FE_OFN1519_acc_fft_data_in_19_), 
	.A0(FE_OFN226_n4525));
   AO22XLTS U2314 (.Y(n6455), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[14] ), 
	.B0(FE_OFN432_n4712), 
	.A1(FE_OFN1727_acc_fir_data_in_14_), 
	.A0(FE_OFN569_n4711));
   AO22XLTS U2309 (.Y(n6450), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[19] ), 
	.B0(FE_OFN424_n4712), 
	.A1(FE_OFN1699_acc_fir_data_in_19_), 
	.A0(FE_OFN562_n4711));
   AO22XLTS U1689 (.Y(n5932), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[8] ), 
	.B0(FE_OFN92_n4526), 
	.A1(FE_OFN1574_acc_fft_data_in_8_), 
	.A0(FE_OFN230_n4525));
   AO22XLTS U1685 (.Y(n5928), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[12] ), 
	.B0(FE_OFN94_n4526), 
	.A1(FE_OFN1555_acc_fft_data_in_12_), 
	.A0(FE_OFN231_n4525));
   AO22XLTS U1679 (.Y(n5922), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[18] ), 
	.B0(FE_OFN85_n4526), 
	.A1(FE_OFN1525_acc_fft_data_in_18_), 
	.A0(FE_OFN226_n4525));
   AO22XLTS U2315 (.Y(n6456), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[13] ), 
	.B0(FE_OFN428_n4712), 
	.A1(FE_OFN1733_acc_fir_data_in_13_), 
	.A0(FE_OFN565_n4711));
   AO22XLTS U1686 (.Y(n5929), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[11] ), 
	.B0(FE_OFN92_n4526), 
	.A1(FE_OFN1559_acc_fft_data_in_11_), 
	.A0(FE_OFN229_n4525));
   AO22XLTS U2313 (.Y(n6454), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[15] ), 
	.B0(FE_OFN429_n4712), 
	.A1(FE_OFN1721_acc_fir_data_in_15_), 
	.A0(FE_OFN566_n4711));
   AO22XLTS U2320 (.Y(n6461), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[8] ), 
	.B0(FE_OFN429_n4712), 
	.A1(FE_OFN1760_acc_fir_data_in_8_), 
	.A0(FE_OFN566_n4711));
   AO22XLTS U2319 (.Y(n6460), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[9] ), 
	.B0(FE_OFN428_n4712), 
	.A1(FE_OFN1752_acc_fir_data_in_9_), 
	.A0(FE_OFN565_n4711));
   AO22XLTS U1690 (.Y(n5933), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[7] ), 
	.B0(FE_OFN86_n4526), 
	.A1(FE_OFN1582_acc_fft_data_in_7_), 
	.A0(FE_OFN223_n4525));
   AO22XLTS U2307 (.Y(n6448), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[21] ), 
	.B0(FE_OFN432_n4712), 
	.A1(FE_OFN1685_acc_fir_data_in_21_), 
	.A0(FE_OFN569_n4711));
   AO22XLTS U2317 (.Y(n6458), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[11] ), 
	.B0(FE_OFN428_n4712), 
	.A1(FE_OFN1742_acc_fir_data_in_11_), 
	.A0(FE_OFN565_n4711));
   AO22XLTS U1684 (.Y(n5927), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[13] ), 
	.B0(FE_OFN93_n4526), 
	.A1(FE_OFN1549_acc_fft_data_in_13_), 
	.A0(FE_OFN230_n4525));
   AO22XLTS U2312 (.Y(n6453), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[16] ), 
	.B0(FE_OFN426_n4712), 
	.A1(FE_OFN1713_acc_fir_data_in_16_), 
	.A0(FE_OFN563_n4711));
   AO22XLTS U1683 (.Y(n5926), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[14] ), 
	.B0(FE_OFN94_n4526), 
	.A1(FE_OFN1546_acc_fft_data_in_14_), 
	.A0(FE_OFN231_n4525));
   AO22XLTS U2308 (.Y(n6449), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[20] ), 
	.B0(n4712), 
	.A1(FE_OFN1692_acc_fir_data_in_20_), 
	.A0(FE_OFN560_n4711));
   AO22XLTS U2316 (.Y(n6457), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[12] ), 
	.B0(FE_OFN432_n4712), 
	.A1(FE_OFN1736_acc_fir_data_in_12_), 
	.A0(FE_OFN569_n4711));
   AO22XLTS U1691 (.Y(n5934), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[6] ), 
	.B0(FE_OFN87_n4526), 
	.A1(FE_OFN1588_acc_fft_data_in_6_), 
	.A0(FE_OFN225_n4525));
   AO22XLTS U2318 (.Y(n6459), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[10] ), 
	.B0(FE_OFN429_n4712), 
	.A1(FE_OFN1748_acc_fir_data_in_10_), 
	.A0(FE_OFN566_n4711));
   AO22XLTS U2306 (.Y(n6447), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[22] ), 
	.B0(FE_OFN432_n4712), 
	.A1(FE_OFN1678_acc_fir_data_in_22_), 
	.A0(FE_OFN569_n4711));
   AO22XLTS U1682 (.Y(n5925), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[15] ), 
	.B0(FE_OFN94_n4526), 
	.A1(FE_OFN1539_acc_fft_data_in_15_), 
	.A0(FE_OFN231_n4525));
   AO22XLTS U1692 (.Y(n5935), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[5] ), 
	.B0(FE_OFN84_n4526), 
	.A1(FE_OFN1593_acc_fft_data_in_5_), 
	.A0(FE_OFN225_n4525));
   AO22XLTS U2305 (.Y(n6446), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[23] ), 
	.B0(FE_OFN424_n4712), 
	.A1(FE_OFN1671_acc_fir_data_in_23_), 
	.A0(FE_OFN563_n4711));
   AO22XLTS U2303 (.Y(n6444), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[25] ), 
	.B0(FE_OFN431_n4712), 
	.A1(FE_OFN1661_acc_fir_data_in_25_), 
	.A0(FE_OFN568_n4711));
   AO22XLTS U1681 (.Y(n5924), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[16] ), 
	.B0(FE_OFN85_n4526), 
	.A1(FE_OFN1537_acc_fft_data_in_16_), 
	.A0(FE_OFN226_n4525));
   AO22XLTS U2302 (.Y(n6443), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[26] ), 
	.B0(FE_OFN431_n4712), 
	.A1(FE_OFN1656_acc_fir_data_in_26_), 
	.A0(FE_OFN568_n4711));
   AO22XLTS U1693 (.Y(n5936), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[4] ), 
	.B0(FE_OFN84_n4526), 
	.A1(FE_OFN1601_acc_fft_data_in_4_), 
	.A0(FE_OFN226_n4525));
   AO22XLTS U1680 (.Y(n5923), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[17] ), 
	.B0(FE_OFN94_n4526), 
	.A1(FE_OFN1529_acc_fft_data_in_17_), 
	.A0(FE_OFN231_n4525));
   AO22XLTS U1670 (.Y(n5913), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[27] ), 
	.B0(FE_OFN89_n4526), 
	.A1(FE_OFN1476_acc_fft_data_in_27_), 
	.A0(FE_OFN224_n4525));
   AO22XLTS U1694 (.Y(n5937), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[3] ), 
	.B0(FE_OFN89_n4526), 
	.A1(FE_OFN1607_acc_fft_data_in_3_), 
	.A0(FE_OFN224_n4525));
   AO22XLTS U1695 (.Y(n5938), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[2] ), 
	.B0(FE_OFN88_n4526), 
	.A1(FE_OFN1614_acc_fft_data_in_2_), 
	.A0(FE_OFN222_n4525));
   AO22XLTS U2304 (.Y(n6445), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[24] ), 
	.B0(FE_OFN431_n4712), 
	.A1(FE_OFN1666_acc_fir_data_in_24_), 
	.A0(FE_OFN568_n4711));
   AO22XLTS U1673 (.Y(n5916), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[24] ), 
	.B0(FE_OFN88_n4526), 
	.A1(FE_OFN1492_acc_fft_data_in_24_), 
	.A0(FE_OFN221_n4525));
   AO22XLTS U1671 (.Y(n5914), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[26] ), 
	.B0(FE_OFN89_n4526), 
	.A1(FE_OFN1481_acc_fft_data_in_26_), 
	.A0(FE_OFN224_n4525));
   AO22XLTS U1696 (.Y(n5939), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[1] ), 
	.B0(FE_OFN86_n4526), 
	.A1(FE_OFN1621_acc_fft_data_in_1_), 
	.A0(FE_OFN222_n4525));
   AO22XLTS U1697 (.Y(n5940), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[0] ), 
	.B0(FE_OFN89_n4526), 
	.A1(FE_OFN1625_acc_fft_data_in_0_), 
	.A0(FE_OFN224_n4525));
   AO22XLTS U1688 (.Y(n5931), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[9] ), 
	.B0(FE_OFN92_n4526), 
	.A1(FE_OFN1569_acc_fft_data_in_9_), 
	.A0(FE_OFN229_n4525));
   AO22XLTS U2301 (.Y(n6442), 
	.B1(\fifo_from_fir/fifo_cell9/sr_out[27] ), 
	.B0(FE_OFN431_n4712), 
	.A1(FE_OFN1653_acc_fir_data_in_27_), 
	.A0(FE_OFN564_n4711));
   AO22XLTS U1672 (.Y(n5915), 
	.B1(\fifo_from_fft/fifo_cell9/sr_out[25] ), 
	.B0(FE_OFN88_n4526), 
	.A1(FE_OFN1485_acc_fft_data_in_25_), 
	.A0(FE_OFN221_n4525));
   OAI21XLTS U2295 (.Y(n4707), 
	.B0(FE_OFN546_n4705), 
	.A1(n4710), 
	.A0(n7554));
   NAND3XLTS U1042 (.Y(n4053), 
	.C(n4139), 
	.B(n4054), 
	.A(n4067));
   NAND3XLTS U898 (.Y(n3878), 
	.C(n3964), 
	.B(n3879), 
	.A(n3892));
   OAI21XLTS U1664 (.Y(n4521), 
	.B0(FE_OFN209_n4519), 
	.A1(n4524), 
	.A0(n7480));
   AO22XLTS U2269 (.Y(n6413), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[22] ), 
	.B0(FE_OFN439_n4706), 
	.A1(FE_OFN1681_acc_fir_data_in_22_), 
	.A0(FE_OFN554_n4705));
   NAND3XLTS U2664 (.Y(n4663), 
	.C(n4799), 
	.B(n4664), 
	.A(FE_OFN546_n4705));
   AOI21X1TS U2293 (.Y(n6436), 
	.B0(FE_OFN803_n7619), 
	.A1(n4707), 
	.A0(\fifo_from_fir/fifo_cell10/controller/valid_read ));
   OAI211XLTS U1043 (.Y(n4138), 
	.C0(n9476), 
	.B0(\fifo_to_fir/hang[13] ), 
	.A1(n4140), 
	.A0(n8787));
   OAI211XLTS U899 (.Y(n3963), 
	.C0(n9480), 
	.B0(\fifo_to_fft/hang[13] ), 
	.A1(n3965), 
	.A0(n8808));
   OAI21XLTS U2294 (.Y(n6437), 
	.B0(n4707), 
	.A1(n4709), 
	.A0(\fifo_from_fir/fifo_cell10/data_out/N35 ));
   AO22XLTS U2270 (.Y(n6414), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[21] ), 
	.B0(FE_OFN436_n4706), 
	.A1(FE_OFN1687_acc_fir_data_in_21_), 
	.A0(FE_OFN550_n4705));
   INVX1TS U3327 (.Y(n4056), 
	.A(n4062));
   NAND3XLTS U2033 (.Y(n4477), 
	.C(n4613), 
	.B(n4478), 
	.A(n4519));
   AO22XLTS U2262 (.Y(n6406), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[29] ), 
	.B0(FE_OFN442_n4706), 
	.A1(FE_OFN1645_acc_fir_data_in_29_), 
	.A0(FE_OFN557_n4705));
   AO22XLTS U1638 (.Y(n5884), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[22] ), 
	.B0(FE_OFN103_n4520), 
	.A1(FE_OFN1501_acc_fft_data_in_22_), 
	.A0(FE_OFN219_n4519));
   OAI21XLTS U1663 (.Y(n5908), 
	.B0(n4521), 
	.A1(n4523), 
	.A0(\fifo_from_fft/fifo_cell10/data_out/N35 ));
   INVX1TS U3470 (.Y(n3881), 
	.A(n3887));
   OAI211XLTS U2665 (.Y(n4798), 
	.C0(n9468), 
	.B0(\fifo_from_fir/hang[9] ), 
	.A1(n4800), 
	.A0(n8875));
   AO22XLTS U2261 (.Y(n6405), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[30] ), 
	.B0(FE_OFN442_n4706), 
	.A1(FE_OFN1637_acc_fir_data_in_30_), 
	.A0(FE_OFN557_n4705));
   AO22XLTS U2271 (.Y(n6415), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[20] ), 
	.B0(FE_OFN433_n4706), 
	.A1(FE_OFN1690_acc_fir_data_in_20_), 
	.A0(FE_OFN549_n4705));
   AO22XLTS U2268 (.Y(n6412), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[23] ), 
	.B0(FE_OFN436_n4706), 
	.A1(FE_OFN1676_acc_fir_data_in_23_), 
	.A0(FE_OFN550_n4705));
   AO22XLTS U1639 (.Y(n5885), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[21] ), 
	.B0(FE_OFN103_n4520), 
	.A1(FE_OFN1507_acc_fft_data_in_21_), 
	.A0(FE_OFN219_n4519));
   AO22XLTS U2260 (.Y(n6404), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[31] ), 
	.B0(FE_OFN442_n4706), 
	.A1(FE_OFN1632_acc_fir_data_in_31_), 
	.A0(FE_OFN557_n4705));
   AOI21X1TS U1662 (.Y(n5907), 
	.B0(FE_OFN820_n7619), 
	.A1(n4521), 
	.A0(\fifo_from_fft/fifo_cell10/controller/valid_read ));
   AO22XLTS U1631 (.Y(n5877), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[29] ), 
	.B0(FE_OFN102_n4520), 
	.A1(FE_OFN1464_acc_fft_data_in_29_), 
	.A0(FE_OFN216_n4519));
   AO22XLTS U2263 (.Y(n6407), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[28] ), 
	.B0(FE_OFN442_n4706), 
	.A1(FE_OFN1650_acc_fir_data_in_28_), 
	.A0(FE_OFN557_n4705));
   AO22XLTS U1637 (.Y(n5883), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[23] ), 
	.B0(FE_OFN97_n4520), 
	.A1(FE_OFN1496_acc_fft_data_in_23_), 
	.A0(FE_OFN213_n4519));
   AO22XLTS U1630 (.Y(n5876), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[30] ), 
	.B0(FE_OFN102_n4520), 
	.A1(FE_OFN1461_acc_fft_data_in_30_), 
	.A0(FE_OFN216_n4519));
   AO22XLTS U1629 (.Y(n5875), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[31] ), 
	.B0(FE_OFN102_n4520), 
	.A1(FE_OFN1455_acc_fft_data_in_31_), 
	.A0(FE_OFN216_n4519));
   AO22XLTS U2274 (.Y(n6418), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[17] ), 
	.B0(FE_OFN435_n4706), 
	.A1(FE_OFN1711_acc_fir_data_in_17_), 
	.A0(FE_OFN551_n4705));
   AO22XLTS U1640 (.Y(n5886), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[20] ), 
	.B0(FE_OFN101_n4520), 
	.A1(FE_OFN1511_acc_fft_data_in_20_), 
	.A0(FE_OFN218_n4519));
   AO22XLTS U2273 (.Y(n6417), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[18] ), 
	.B0(FE_OFN435_n4706), 
	.A1(FE_OFN1703_acc_fir_data_in_18_), 
	.A0(FE_OFN551_n4705));
   OAI211XLTS U2034 (.Y(n4612), 
	.C0(n9471), 
	.B0(\fifo_from_fft/hang[9] ), 
	.A1(n4614), 
	.A0(n8842));
   AO22XLTS U2275 (.Y(n6419), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[16] ), 
	.B0(FE_OFN435_n4706), 
	.A1(FE_OFN1712_acc_fir_data_in_16_), 
	.A0(FE_OFN551_n4705));
   AO22XLTS U2272 (.Y(n6416), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[19] ), 
	.B0(FE_OFN433_n4706), 
	.A1(FE_OFN1701_acc_fir_data_in_19_), 
	.A0(FE_OFN549_n4705));
   AO22XLTS U2280 (.Y(n6424), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[11] ), 
	.B0(FE_OFN440_n4706), 
	.A1(FE_OFN1745_acc_fir_data_in_11_), 
	.A0(FE_OFN556_n4705));
   AO22XLTS U1641 (.Y(n5887), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[19] ), 
	.B0(FE_OFN98_n4520), 
	.A1(FE_OFN1519_acc_fft_data_in_19_), 
	.A0(FE_OFN215_n4519));
   AO22XLTS U1632 (.Y(n5878), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[28] ), 
	.B0(FE_OFN103_n4520), 
	.A1(FE_OFN1472_acc_fft_data_in_28_), 
	.A0(FE_OFN219_n4519));
   AO22XLTS U2277 (.Y(n6421), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[14] ), 
	.B0(FE_OFN436_n4706), 
	.A1(FE_OFN1728_acc_fir_data_in_14_), 
	.A0(FE_OFN550_n4705));
   AO22XLTS U2283 (.Y(n6427), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[8] ), 
	.B0(FE_OFN440_n4706), 
	.A1(FE_OFN1757_acc_fir_data_in_8_), 
	.A0(FE_OFN556_n4705));
   AO22XLTS U2284 (.Y(n6428), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[7] ), 
	.B0(FE_OFN437_n4706), 
	.A1(FE_OFN1763_acc_fir_data_in_7_), 
	.A0(FE_OFN553_n4705));
   AO22XLTS U2286 (.Y(n6430), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[5] ), 
	.B0(FE_OFN438_n4706), 
	.A1(FE_OFN1782_acc_fir_data_in_5_), 
	.A0(FE_OFN552_n4705));
   AO22XLTS U2291 (.Y(n6435), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[0] ), 
	.B0(FE_OFN437_n4706), 
	.A1(FE_OFN1810_acc_fir_data_in_0_), 
	.A0(FE_OFN553_n4705));
   AO22XLTS U1644 (.Y(n5890), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[16] ), 
	.B0(FE_OFN100_n4520), 
	.A1(FE_OFN1536_acc_fft_data_in_16_), 
	.A0(FE_OFN217_n4519));
   AO22XLTS U2285 (.Y(n6429), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[6] ), 
	.B0(FE_OFN434_n4706), 
	.A1(FE_OFN1770_acc_fir_data_in_6_), 
	.A0(FE_OFN548_n4705));
   AO22XLTS U2266 (.Y(n6410), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[25] ), 
	.B0(FE_OFN441_n4706), 
	.A1(FE_OFN1665_acc_fir_data_in_25_), 
	.A0(FE_OFN555_n4705));
   AO22XLTS U2290 (.Y(n6434), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[1] ), 
	.B0(n4706), 
	.A1(FE_OFN1807_acc_fir_data_in_1_), 
	.A0(n4705));
   AO22XLTS U2288 (.Y(n6432), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[3] ), 
	.B0(n4706), 
	.A1(FE_OFN1794_acc_fir_data_in_3_), 
	.A0(FE_OFN547_n4705));
   AO22XLTS U2287 (.Y(n6431), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[4] ), 
	.B0(FE_OFN434_n4706), 
	.A1(FE_OFN1788_acc_fir_data_in_4_), 
	.A0(FE_OFN548_n4705));
   AO22XLTS U1643 (.Y(n5889), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[17] ), 
	.B0(FE_OFN100_n4520), 
	.A1(FE_OFN1531_acc_fft_data_in_17_), 
	.A0(FE_OFN217_n4519));
   AO22XLTS U2289 (.Y(n6433), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[2] ), 
	.B0(FE_OFN437_n4706), 
	.A1(FE_OFN1795_acc_fir_data_in_2_), 
	.A0(FE_OFN553_n4705));
   AO22XLTS U2279 (.Y(n6423), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[12] ), 
	.B0(FE_OFN439_n4706), 
	.A1(FE_OFN1736_acc_fir_data_in_12_), 
	.A0(FE_OFN554_n4705));
   AO22XLTS U2278 (.Y(n6422), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[13] ), 
	.B0(FE_OFN440_n4706), 
	.A1(FE_OFN1731_acc_fir_data_in_13_), 
	.A0(FE_OFN556_n4705));
   AO22XLTS U2265 (.Y(n6409), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[26] ), 
	.B0(FE_OFN441_n4706), 
	.A1(FE_OFN1658_acc_fir_data_in_26_), 
	.A0(FE_OFN555_n4705));
   AO22XLTS U2267 (.Y(n6411), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[24] ), 
	.B0(FE_OFN441_n4706), 
	.A1(FE_OFN1670_acc_fir_data_in_24_), 
	.A0(FE_OFN555_n4705));
   AO22XLTS U1642 (.Y(n5888), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[18] ), 
	.B0(FE_OFN101_n4520), 
	.A1(FE_OFN1522_acc_fft_data_in_18_), 
	.A0(FE_OFN218_n4519));
   AO22XLTS U2282 (.Y(n6426), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[9] ), 
	.B0(FE_OFN440_n4706), 
	.A1(FE_OFN1751_acc_fir_data_in_9_), 
	.A0(FE_OFN556_n4705));
   AO22XLTS U2264 (.Y(n6408), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[27] ), 
	.B0(FE_OFN438_n4706), 
	.A1(FE_OFN1655_acc_fir_data_in_27_), 
	.A0(FE_OFN552_n4705));
   AO22XLTS U2276 (.Y(n6420), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[15] ), 
	.B0(FE_OFN439_n4706), 
	.A1(FE_OFN1719_acc_fir_data_in_15_), 
	.A0(FE_OFN554_n4705));
   AO22XLTS U2281 (.Y(n6425), 
	.B1(\fifo_from_fir/fifo_cell10/sr_out[10] ), 
	.B0(FE_OFN439_n4706), 
	.A1(FE_OFN1746_acc_fir_data_in_10_), 
	.A0(FE_OFN554_n4705));
   AO22XLTS U1649 (.Y(n5895), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[11] ), 
	.B0(FE_OFN104_n4520), 
	.A1(FE_OFN1561_acc_fft_data_in_11_), 
	.A0(FE_OFN220_n4519));
   AO22XLTS U1646 (.Y(n5892), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[14] ), 
	.B0(FE_OFN98_n4520), 
	.A1(FE_OFN1547_acc_fft_data_in_14_), 
	.A0(FE_OFN215_n4519));
   AO22XLTS U1635 (.Y(n5881), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[25] ), 
	.B0(n4520), 
	.A1(FE_OFN1487_acc_fft_data_in_25_), 
	.A0(FE_OFN210_n4519));
   AO22XLTS U1647 (.Y(n5893), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[13] ), 
	.B0(FE_OFN101_n4520), 
	.A1(FE_OFN1552_acc_fft_data_in_13_), 
	.A0(FE_OFN218_n4519));
   AO22XLTS U1653 (.Y(n5899), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[7] ), 
	.B0(FE_OFN97_n4520), 
	.A1(FE_OFN1583_acc_fft_data_in_7_), 
	.A0(FE_OFN212_n4519));
   OAI21XLTS U2258 (.Y(n4701), 
	.B0(FE_OFN534_n4699), 
	.A1(n4704), 
	.A0(n7549));
   AO22XLTS U1659 (.Y(n5905), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[1] ), 
	.B0(FE_OFN96_n4520), 
	.A1(FE_OFN1620_acc_fft_data_in_1_), 
	.A0(FE_OFN211_n4519));
   AO22XLTS U1633 (.Y(n5879), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[27] ), 
	.B0(FE_OFN96_n4520), 
	.A1(FE_OFN1477_acc_fft_data_in_27_), 
	.A0(FE_OFN211_n4519));
   AO22XLTS U1645 (.Y(n5891), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[15] ), 
	.B0(FE_OFN101_n4520), 
	.A1(FE_OFN1541_acc_fft_data_in_15_), 
	.A0(FE_OFN218_n4519));
   AO22XLTS U1660 (.Y(n5906), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[0] ), 
	.B0(FE_OFN99_n4520), 
	.A1(FE_OFN1625_acc_fft_data_in_0_), 
	.A0(FE_OFN214_n4519));
   OAI211XLTS U897 (.Y(n3962), 
	.C0(n9480), 
	.B0(\fifo_to_fft/hang[14] ), 
	.A1(n3880), 
	.A0(n8810));
   AO22XLTS U1648 (.Y(n5894), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[12] ), 
	.B0(FE_OFN100_n4520), 
	.A1(FE_OFN1558_acc_fft_data_in_12_), 
	.A0(FE_OFN217_n4519));
   AO22XLTS U1651 (.Y(n5897), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[9] ), 
	.B0(FE_OFN104_n4520), 
	.A1(FE_OFN1573_acc_fft_data_in_9_), 
	.A0(FE_OFN220_n4519));
   AO22XLTS U1650 (.Y(n5896), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[10] ), 
	.B0(FE_OFN104_n4520), 
	.A1(FE_OFN1568_acc_fft_data_in_10_), 
	.A0(FE_OFN220_n4519));
   AO22XLTS U1634 (.Y(n5880), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[26] ), 
	.B0(FE_OFN99_n4520), 
	.A1(FE_OFN1482_acc_fft_data_in_26_), 
	.A0(FE_OFN214_n4519));
   AO22XLTS U1656 (.Y(n5902), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[4] ), 
	.B0(FE_OFN95_n4520), 
	.A1(FE_OFN1599_acc_fft_data_in_4_), 
	.A0(FE_OFN213_n4519));
   AO22XLTS U1654 (.Y(n5900), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[6] ), 
	.B0(FE_OFN97_n4520), 
	.A1(FE_OFN1587_acc_fft_data_in_6_), 
	.A0(FE_OFN213_n4519));
   AO22XLTS U1636 (.Y(n5882), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[24] ), 
	.B0(n4520), 
	.A1(FE_OFN1491_acc_fft_data_in_24_), 
	.A0(n4519));
   AO22XLTS U1652 (.Y(n5898), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[8] ), 
	.B0(FE_OFN104_n4520), 
	.A1(FE_OFN1578_acc_fft_data_in_8_), 
	.A0(FE_OFN220_n4519));
   AO22XLTS U1657 (.Y(n5903), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[3] ), 
	.B0(FE_OFN99_n4520), 
	.A1(FE_OFN1607_acc_fft_data_in_3_), 
	.A0(FE_OFN214_n4519));
   AO22XLTS U1658 (.Y(n5904), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[2] ), 
	.B0(FE_OFN96_n4520), 
	.A1(FE_OFN1614_acc_fft_data_in_2_), 
	.A0(FE_OFN211_n4519));
   AO22XLTS U1655 (.Y(n5901), 
	.B1(\fifo_from_fft/fifo_cell10/sr_out[5] ), 
	.B0(FE_OFN97_n4520), 
	.A1(FE_OFN1593_acc_fft_data_in_5_), 
	.A0(FE_OFN212_n4519));
   AOI21X1TS U2256 (.Y(n6402), 
	.B0(FE_OFN808_n7619), 
	.A1(n4701), 
	.A0(\fifo_from_fir/fifo_cell11/controller/valid_read ));
   NAND3XLTS U2662 (.Y(n4665), 
	.C(n4796), 
	.B(n4666), 
	.A(FE_OFN534_n4699));
   OAI21XLTS U1627 (.Y(n4515), 
	.B0(FE_OFN199_n4513), 
	.A1(n4518), 
	.A0(n7475));
   OAI31XLTS U896 (.Y(n5516), 
	.B0(n3962), 
	.A2(n3880), 
	.A1(n3881), 
	.A0(\fifo_to_fft/hang[14] ));
   OAI31XLTS U1040 (.Y(n5568), 
	.B0(n4137), 
	.A2(n4055), 
	.A1(n4056), 
	.A0(\fifo_to_fir/hang[14] ));
   OAI21XLTS U2257 (.Y(n6403), 
	.B0(n4701), 
	.A1(n4703), 
	.A0(\fifo_from_fir/fifo_cell11/data_out/N35 ));
   AO22XLTS U2242 (.Y(n6389), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[12] ), 
	.B0(FE_OFN532_n4700), 
	.A1(FE_OFN1739_acc_fir_data_in_12_), 
	.A0(FE_OFN544_n4699));
   OAI211XLTS U2663 (.Y(n4795), 
	.C0(n9468), 
	.B0(\fifo_from_fir/hang[10] ), 
	.A1(n4797), 
	.A0(n8874));
   AO22XLTS U2223 (.Y(n6370), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[31] ), 
	.B0(FE_OFN533_n4700), 
	.A1(FE_OFN1629_acc_fir_data_in_31_), 
	.A0(FE_OFN545_n4699));
   AOI21X1TS U1625 (.Y(n5873), 
	.B0(FE_OFN820_n7619), 
	.A1(n4515), 
	.A0(\fifo_from_fft/fifo_cell11/controller/valid_read ));
   AO22XLTS U2240 (.Y(n6387), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[14] ), 
	.B0(FE_OFN532_n4700), 
	.A1(FE_OFN1730_acc_fir_data_in_14_), 
	.A0(FE_OFN544_n4699));
   NAND3XLTS U2031 (.Y(n4479), 
	.C(n4610), 
	.B(n4480), 
	.A(FE_OFN199_n4513));
   AO22XLTS U2226 (.Y(n6373), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[28] ), 
	.B0(FE_OFN533_n4700), 
	.A1(FE_OFN1649_acc_fir_data_in_28_), 
	.A0(FE_OFN545_n4699));
   OAI21XLTS U1626 (.Y(n5874), 
	.B0(n4515), 
	.A1(n4517), 
	.A0(\fifo_from_fft/fifo_cell11/data_out/N35 ));
   AO22XLTS U2225 (.Y(n6372), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[29] ), 
	.B0(FE_OFN533_n4700), 
	.A1(FE_OFN1644_acc_fir_data_in_29_), 
	.A0(FE_OFN545_n4699));
   AO22XLTS U2224 (.Y(n6371), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[30] ), 
	.B0(FE_OFN533_n4700), 
	.A1(FE_OFN1636_acc_fir_data_in_30_), 
	.A0(FE_OFN545_n4699));
   AO22XLTS U2241 (.Y(n6388), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[13] ), 
	.B0(FE_OFN528_n4700), 
	.A1(FE_OFN1733_acc_fir_data_in_13_), 
	.A0(FE_OFN539_n4699));
   AO22XLTS U2239 (.Y(n6386), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[15] ), 
	.B0(FE_OFN532_n4700), 
	.A1(FE_OFN1723_acc_fir_data_in_15_), 
	.A0(FE_OFN544_n4699));
   AO22XLTS U1595 (.Y(n5844), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[28] ), 
	.B0(FE_OFN195_n4514), 
	.A1(FE_OFN1472_acc_fft_data_in_28_), 
	.A0(FE_OFN207_n4513));
   AO22XLTS U1593 (.Y(n5842), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[30] ), 
	.B0(FE_OFN192_n4514), 
	.A1(FE_OFN1461_acc_fft_data_in_30_), 
	.A0(FE_OFN204_n4513));
   AO22XLTS U2234 (.Y(n6381), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[20] ), 
	.B0(FE_OFN525_n4700), 
	.A1(FE_OFN1693_acc_fir_data_in_20_), 
	.A0(FE_OFN538_n4699));
   AO22XLTS U2252 (.Y(n6399), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[2] ), 
	.B0(FE_OFN524_n4700), 
	.A1(FE_OFN1800_acc_fir_data_in_2_), 
	.A0(FE_OFN537_n4699));
   AOI21X1TS U778 (.Y(n5454), 
	.B0(FE_OFN798_n7619), 
	.A1(n3808), 
	.A0(\fifo_to_fir/fifo_cell0/controller/valid_read ));
   AO22XLTS U2237 (.Y(n6384), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[17] ), 
	.B0(FE_OFN523_n4700), 
	.A1(FE_OFN1709_acc_fir_data_in_17_), 
	.A0(FE_OFN536_n4699));
   AO22XLTS U2250 (.Y(n6397), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[4] ), 
	.B0(FE_OFN526_n4700), 
	.A1(FE_OFN1786_acc_fir_data_in_4_), 
	.A0(FE_OFN537_n4699));
   AO22XLTS U2238 (.Y(n6385), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[16] ), 
	.B0(FE_OFN527_n4700), 
	.A1(FE_OFN1718_acc_fir_data_in_16_), 
	.A0(FE_OFN536_n4699));
   AO22XLTS U2249 (.Y(n6396), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[5] ), 
	.B0(FE_OFN529_n4700), 
	.A1(FE_OFN1781_acc_fir_data_in_5_), 
	.A0(FE_OFN540_n4699));
   AO22XLTS U2246 (.Y(n6393), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[8] ), 
	.B0(FE_OFN530_n4700), 
	.A1(FE_OFN1761_acc_fir_data_in_8_), 
	.A0(FE_OFN542_n4699));
   AO22XLTS U2227 (.Y(n6374), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[27] ), 
	.B0(FE_OFN531_n4700), 
	.A1(FE_OFN1654_acc_fir_data_in_27_), 
	.A0(FE_OFN541_n4699));
   AO22XLTS U2228 (.Y(n6375), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[26] ), 
	.B0(FE_OFN531_n4700), 
	.A1(FE_OFN1660_acc_fir_data_in_26_), 
	.A0(FE_OFN541_n4699));
   AO22XLTS U2229 (.Y(n6376), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[25] ), 
	.B0(FE_OFN529_n4700), 
	.A1(FE_OFN1663_acc_fir_data_in_25_), 
	.A0(FE_OFN543_n4699));
   AO22XLTS U2253 (.Y(n6400), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[1] ), 
	.B0(n4700), 
	.A1(FE_OFN1807_acc_fir_data_in_1_), 
	.A0(n4699));
   AO22XLTS U2230 (.Y(n6377), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[24] ), 
	.B0(FE_OFN529_n4700), 
	.A1(FE_OFN1668_acc_fir_data_in_24_), 
	.A0(FE_OFN543_n4699));
   AO22XLTS U2254 (.Y(n6401), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[0] ), 
	.B0(FE_OFN524_n4700), 
	.A1(FE_OFN1811_acc_fir_data_in_0_), 
	.A0(FE_OFN537_n4699));
   AO22XLTS U2245 (.Y(n6392), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[9] ), 
	.B0(FE_OFN530_n4700), 
	.A1(FE_OFN1754_acc_fir_data_in_9_), 
	.A0(FE_OFN542_n4699));
   AO22XLTS U2231 (.Y(n6378), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[23] ), 
	.B0(FE_OFN525_n4700), 
	.A1(FE_OFN1673_acc_fir_data_in_23_), 
	.A0(FE_OFN538_n4699));
   OAI211XLTS U2032 (.Y(n4609), 
	.C0(n9472), 
	.B0(\fifo_from_fft/hang[10] ), 
	.A1(n4611), 
	.A0(n8841));
   AO22XLTS U2232 (.Y(n6379), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[22] ), 
	.B0(FE_OFN532_n4700), 
	.A1(FE_OFN1681_acc_fir_data_in_22_), 
	.A0(FE_OFN544_n4699));
   AO22XLTS U2251 (.Y(n6398), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[3] ), 
	.B0(FE_OFN524_n4700), 
	.A1(FE_OFN1790_acc_fir_data_in_3_), 
	.A0(FE_OFN535_n4699));
   AO22XLTS U2247 (.Y(n6394), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[7] ), 
	.B0(FE_OFN526_n4700), 
	.A1(FE_OFN1765_acc_fir_data_in_7_), 
	.A0(FE_OFN540_n4699));
   AO22XLTS U1610 (.Y(n5859), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[13] ), 
	.B0(FE_OFN194_n4514), 
	.A1(FE_OFN1551_acc_fft_data_in_13_), 
	.A0(FE_OFN206_n4513));
   AO22XLTS U2233 (.Y(n6380), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[21] ), 
	.B0(FE_OFN527_n4700), 
	.A1(FE_OFN1689_acc_fir_data_in_21_), 
	.A0(FE_OFN538_n4699));
   AO22XLTS U1592 (.Y(n5841), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[31] ), 
	.B0(FE_OFN192_n4514), 
	.A1(FE_OFN1457_acc_fft_data_in_31_), 
	.A0(FE_OFN204_n4513));
   AO22XLTS U2243 (.Y(n6390), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[11] ), 
	.B0(FE_OFN528_n4700), 
	.A1(FE_OFN1744_acc_fir_data_in_11_), 
	.A0(FE_OFN539_n4699));
   AO22XLTS U2236 (.Y(n6383), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[18] ), 
	.B0(FE_OFN527_n4700), 
	.A1(FE_OFN1705_acc_fir_data_in_18_), 
	.A0(FE_OFN539_n4699));
   AO22XLTS U2248 (.Y(n6395), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[6] ), 
	.B0(FE_OFN526_n4700), 
	.A1(FE_OFN1776_acc_fir_data_in_6_), 
	.A0(FE_OFN540_n4699));
   AO22XLTS U2235 (.Y(n6382), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[19] ), 
	.B0(FE_OFN523_n4700), 
	.A1(FE_OFN1700_acc_fir_data_in_19_), 
	.A0(FE_OFN535_n4699));
   AO22XLTS U2244 (.Y(n6391), 
	.B1(\fifo_from_fir/fifo_cell11/sr_out[10] ), 
	.B0(FE_OFN530_n4700), 
	.A1(FE_OFN1749_acc_fir_data_in_10_), 
	.A0(FE_OFN542_n4699));
   AO22XLTS U1608 (.Y(n5857), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[15] ), 
	.B0(FE_OFN194_n4514), 
	.A1(FE_OFN1540_acc_fft_data_in_15_), 
	.A0(FE_OFN206_n4513));
   AO22XLTS U1611 (.Y(n5860), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[12] ), 
	.B0(FE_OFN194_n4514), 
	.A1(FE_OFN1556_acc_fft_data_in_12_), 
	.A0(FE_OFN205_n4513));
   AO22XLTS U1609 (.Y(n5858), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[14] ), 
	.B0(FE_OFN194_n4514), 
	.A1(FE_OFN1544_acc_fft_data_in_14_), 
	.A0(FE_OFN206_n4513));
   AO22XLTS U1594 (.Y(n5843), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[29] ), 
	.B0(FE_OFN192_n4514), 
	.A1(FE_OFN1466_acc_fft_data_in_29_), 
	.A0(FE_OFN204_n4513));
   AO22XLTS U1601 (.Y(n5850), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[22] ), 
	.B0(FE_OFN195_n4514), 
	.A1(FE_OFN1501_acc_fft_data_in_22_), 
	.A0(FE_OFN207_n4513));
   AO22XLTS U1622 (.Y(n5871), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[1] ), 
	.B0(FE_OFN189_n4514), 
	.A1(FE_OFN1618_acc_fft_data_in_1_), 
	.A0(FE_OFN200_n4513));
   AO22XLTS U1603 (.Y(n5852), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[20] ), 
	.B0(FE_OFN190_n4514), 
	.A1(FE_OFN1511_acc_fft_data_in_20_), 
	.A0(FE_OFN203_n4513));
   AO22XLTS U1623 (.Y(n5872), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[0] ), 
	.B0(FE_OFN191_n4514), 
	.A1(FE_OFN1624_acc_fft_data_in_0_), 
	.A0(FE_OFN201_n4513));
   AO22XLTS U1604 (.Y(n5853), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[19] ), 
	.B0(FE_OFN193_n4514), 
	.A1(FE_OFN1516_acc_fft_data_in_19_), 
	.A0(FE_OFN205_n4513));
   AO22XLTS U1597 (.Y(n5846), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[26] ), 
	.B0(FE_OFN191_n4514), 
	.A1(FE_OFN1481_acc_fft_data_in_26_), 
	.A0(FE_OFN201_n4513));
   AO22XLTS U1621 (.Y(n5870), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[2] ), 
	.B0(FE_OFN189_n4514), 
	.A1(FE_OFN1612_acc_fft_data_in_2_), 
	.A0(FE_OFN197_n4513));
   AO22XLTS U1615 (.Y(n5864), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[8] ), 
	.B0(FE_OFN196_n4514), 
	.A1(FE_OFN1578_acc_fft_data_in_8_), 
	.A0(FE_OFN208_n4513));
   AO22XLTS U1599 (.Y(n5848), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[24] ), 
	.B0(FE_OFN187_n4514), 
	.A1(FE_OFN1491_acc_fft_data_in_24_), 
	.A0(FE_OFN197_n4513));
   AO22XLTS U1616 (.Y(n5865), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[7] ), 
	.B0(FE_OFN187_n4514), 
	.A1(FE_OFN1584_acc_fft_data_in_7_), 
	.A0(FE_OFN198_n4513));
   AO22XLTS U1600 (.Y(n5849), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[23] ), 
	.B0(FE_OFN190_n4514), 
	.A1(FE_OFN1497_acc_fft_data_in_23_), 
	.A0(FE_OFN202_n4513));
   AO22XLTS U1605 (.Y(n5854), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[18] ), 
	.B0(FE_OFN190_n4514), 
	.A1(FE_OFN1522_acc_fft_data_in_18_), 
	.A0(FE_OFN203_n4513));
   AO22XLTS U1606 (.Y(n5855), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[17] ), 
	.B0(FE_OFN193_n4514), 
	.A1(FE_OFN1531_acc_fft_data_in_17_), 
	.A0(FE_OFN205_n4513));
   AO22XLTS U1612 (.Y(n5861), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[11] ), 
	.B0(FE_OFN196_n4514), 
	.A1(FE_OFN1561_acc_fft_data_in_11_), 
	.A0(FE_OFN208_n4513));
   AO22XLTS U1620 (.Y(n5869), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[3] ), 
	.B0(FE_OFN191_n4514), 
	.A1(FE_OFN1605_acc_fft_data_in_3_), 
	.A0(FE_OFN201_n4513));
   AO22XLTS U1619 (.Y(n5868), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[4] ), 
	.B0(FE_OFN188_n4514), 
	.A1(FE_OFN1601_acc_fft_data_in_4_), 
	.A0(FE_OFN198_n4513));
   AO22XLTS U1602 (.Y(n5851), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[21] ), 
	.B0(FE_OFN195_n4514), 
	.A1(FE_OFN1509_acc_fft_data_in_21_), 
	.A0(FE_OFN207_n4513));
   AO22XLTS U1607 (.Y(n5856), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[16] ), 
	.B0(FE_OFN193_n4514), 
	.A1(FE_OFN1536_acc_fft_data_in_16_), 
	.A0(FE_OFN205_n4513));
   AO22XLTS U1613 (.Y(n5862), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[10] ), 
	.B0(FE_OFN196_n4514), 
	.A1(FE_OFN1568_acc_fft_data_in_10_), 
	.A0(FE_OFN208_n4513));
   AO22XLTS U1598 (.Y(n5847), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[25] ), 
	.B0(FE_OFN187_n4514), 
	.A1(FE_OFN1485_acc_fft_data_in_25_), 
	.A0(FE_OFN197_n4513));
   AO22XLTS U1596 (.Y(n5845), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[27] ), 
	.B0(FE_OFN189_n4514), 
	.A1(FE_OFN1476_acc_fft_data_in_27_), 
	.A0(FE_OFN200_n4513));
   AO22XLTS U1614 (.Y(n5863), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[9] ), 
	.B0(FE_OFN196_n4514), 
	.A1(FE_OFN1573_acc_fft_data_in_9_), 
	.A0(FE_OFN208_n4513));
   AO22XLTS U1617 (.Y(n5866), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[6] ), 
	.B0(FE_OFN188_n4514), 
	.A1(FE_OFN1590_acc_fft_data_in_6_), 
	.A0(FE_OFN202_n4513));
   AO22XLTS U1618 (.Y(n5867), 
	.B1(\fifo_from_fft/fifo_cell11/sr_out[5] ), 
	.B0(FE_OFN188_n4514), 
	.A1(FE_OFN1595_acc_fft_data_in_5_), 
	.A0(FE_OFN202_n4513));
   OAI21XLTS U2221 (.Y(n4695), 
	.B0(n4693), 
	.A1(n4698), 
	.A0(n7544));
   NAND2X1TS U3540 (.Y(\fifo_to_fft/fifo_cell0/reg_ptok/N22 ), 
	.B(n5250), 
	.A(n9514));
   NAND2XLTS U3396 (.Y(\fifo_to_fir/fifo_cell0/reg_ptok/N22 ), 
	.B(n5208), 
	.A(n9515));
   AO22XLTS U2195 (.Y(n6345), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[22] ), 
	.B0(FE_OFN449_n4694), 
	.A1(FE_OFN1678_acc_fir_data_in_22_), 
	.A0(FE_OFN522_n4693));
   OAI21X1TS U1590 (.Y(n4509), 
	.B0(FE_OFN175_n4507), 
	.A1(n4512), 
	.A0(n7470));
   NAND3XLTS U2660 (.Y(n4667), 
	.C(n4793), 
	.B(n4668), 
	.A(FE_OFN511_n4693));
   AO22XLTS U2196 (.Y(n6346), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[21] ), 
	.B0(FE_OFN449_n4694), 
	.A1(FE_OFN1688_acc_fir_data_in_21_), 
	.A0(FE_OFN522_n4693));
   OAI21XLTS U2220 (.Y(n6369), 
	.B0(n4695), 
	.A1(n4697), 
	.A0(\fifo_from_fir/fifo_cell12/data_out/N35 ));
   AO22XLTS U2186 (.Y(n6336), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[31] ), 
	.B0(FE_OFN452_n4694), 
	.A1(FE_OFN1631_acc_fir_data_in_31_), 
	.A0(FE_OFN514_n4693));
   AO22XLTS U2187 (.Y(n6337), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[30] ), 
	.B0(FE_OFN452_n4694), 
	.A1(FE_OFN1635_acc_fir_data_in_30_), 
	.A0(FE_OFN514_n4693));
   OAI211XLTS U2661 (.Y(n4792), 
	.C0(n9465), 
	.B0(\fifo_from_fir/hang[11] ), 
	.A1(n4794), 
	.A0(n8874));
   AO22XLTS U1565 (.Y(n5817), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[21] ), 
	.B0(FE_OFN113_n4508), 
	.A1(FE_OFN1509_acc_fft_data_in_21_), 
	.A0(FE_OFN185_n4507));
   NAND3XLTS U2029 (.Y(n4481), 
	.C(n4607), 
	.B(n4482), 
	.A(FE_OFN175_n4507));
   AO22XLTS U2188 (.Y(n6338), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[29] ), 
	.B0(FE_OFN452_n4694), 
	.A1(FE_OFN1643_acc_fir_data_in_29_), 
	.A0(FE_OFN514_n4693));
   AO22XLTS U2197 (.Y(n6347), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[20] ), 
	.B0(FE_OFN443_n4694), 
	.A1(FE_OFN1693_acc_fir_data_in_20_), 
	.A0(FE_OFN517_n4693));
   AO22XLTS U1564 (.Y(n5816), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[22] ), 
	.B0(FE_OFN113_n4508), 
	.A1(FE_OFN1500_acc_fft_data_in_22_), 
	.A0(FE_OFN185_n4507));
   AO22XLTS U2194 (.Y(n6344), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[23] ), 
	.B0(n4694), 
	.A1(FE_OFN1673_acc_fir_data_in_23_), 
	.A0(FE_OFN518_n4693));
   OAI21XLTS U1589 (.Y(n5840), 
	.B0(n4509), 
	.A1(n4511), 
	.A0(\fifo_from_fft/fifo_cell12/data_out/N35 ));
   AO22XLTS U1566 (.Y(n5818), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[20] ), 
	.B0(FE_OFN110_n4508), 
	.A1(FE_OFN1511_acc_fft_data_in_20_), 
	.A0(FE_OFN181_n4507));
   AO22XLTS U1556 (.Y(n5808), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[30] ), 
	.B0(FE_OFN111_n4508), 
	.A1(FE_OFN1461_acc_fft_data_in_30_), 
	.A0(FE_OFN182_n4507));
   AO22XLTS U2199 (.Y(n6349), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[18] ), 
	.B0(FE_OFN444_n4694), 
	.A1(FE_OFN1706_acc_fir_data_in_18_), 
	.A0(FE_OFN519_n4693));
   AO22XLTS U2198 (.Y(n6348), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[19] ), 
	.B0(FE_OFN443_n4694), 
	.A1(FE_OFN1700_acc_fir_data_in_19_), 
	.A0(FE_OFN517_n4693));
   OAI211XLTS U2030 (.Y(n4606), 
	.C0(n9472), 
	.B0(\fifo_from_fft/hang[11] ), 
	.A1(n4608), 
	.A0(n8841));
   AO22XLTS U1563 (.Y(n5815), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[23] ), 
	.B0(FE_OFN108_n4508), 
	.A1(FE_OFN1494_acc_fft_data_in_23_), 
	.A0(FE_OFN180_n4507));
   AO22XLTS U1557 (.Y(n5809), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[29] ), 
	.B0(FE_OFN111_n4508), 
	.A1(FE_OFN1466_acc_fft_data_in_29_), 
	.A0(FE_OFN184_n4507));
   AO22XLTS U2201 (.Y(n6351), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[16] ), 
	.B0(FE_OFN444_n4694), 
	.A1(FE_OFN1717_acc_fir_data_in_16_), 
	.A0(FE_OFN519_n4693));
   AO22XLTS U2200 (.Y(n6350), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[17] ), 
	.B0(FE_OFN444_n4694), 
	.A1(FE_OFN1710_acc_fir_data_in_17_), 
	.A0(FE_OFN519_n4693));
   AO22XLTS U2189 (.Y(n6339), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[28] ), 
	.B0(FE_OFN452_n4694), 
	.A1(FE_OFN1650_acc_fir_data_in_28_), 
	.A0(FE_OFN514_n4693));
   AO22XLTS U1555 (.Y(n5807), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[31] ), 
	.B0(FE_OFN111_n4508), 
	.A1(FE_OFN1457_acc_fft_data_in_31_), 
	.A0(FE_OFN184_n4507));
   AO22XLTS U2209 (.Y(n6359), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[8] ), 
	.B0(FE_OFN447_n4694), 
	.A1(FE_OFN1760_acc_fir_data_in_8_), 
	.A0(FE_OFN521_n4693));
   AO22XLTS U2214 (.Y(n6364), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[3] ), 
	.B0(FE_OFN445_n4694), 
	.A1(FE_OFN1792_acc_fir_data_in_3_), 
	.A0(FE_OFN516_n4693));
   AO22XLTS U2206 (.Y(n6356), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[11] ), 
	.B0(FE_OFN446_n4694), 
	.A1(FE_OFN1743_acc_fir_data_in_11_), 
	.A0(FE_OFN520_n4693));
   AO22XLTS U2205 (.Y(n6355), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[12] ), 
	.B0(FE_OFN449_n4694), 
	.A1(FE_OFN1738_acc_fir_data_in_12_), 
	.A0(FE_OFN522_n4693));
   AO22XLTS U2217 (.Y(n6367), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[0] ), 
	.B0(FE_OFN445_n4694), 
	.A1(FE_OFN1813_acc_fir_data_in_0_), 
	.A0(FE_OFN516_n4693));
   AO22XLTS U2203 (.Y(n6353), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[14] ), 
	.B0(FE_OFN449_n4694), 
	.A1(FE_OFN1725_acc_fir_data_in_14_), 
	.A0(FE_OFN522_n4693));
   AO22XLTS U1558 (.Y(n5810), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[28] ), 
	.B0(FE_OFN113_n4508), 
	.A1(FE_OFN1470_acc_fft_data_in_28_), 
	.A0(FE_OFN184_n4507));
   AO22XLTS U1567 (.Y(n5819), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[19] ), 
	.B0(FE_OFN108_n4508), 
	.A1(FE_OFN1518_acc_fft_data_in_19_), 
	.A0(FE_OFN180_n4507));
   AO22XLTS U1569 (.Y(n5821), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[17] ), 
	.B0(FE_OFN112_n4508), 
	.A1(FE_OFN1528_acc_fft_data_in_17_), 
	.A0(FE_OFN183_n4507));
   AO22XLTS U2211 (.Y(n6361), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[6] ), 
	.B0(FE_OFN448_n4694), 
	.A1(FE_OFN1771_acc_fir_data_in_6_), 
	.A0(FE_OFN513_n4693));
   AO22XLTS U2216 (.Y(n6366), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[1] ), 
	.B0(FE_OFN443_n4694), 
	.A1(FE_OFN1803_acc_fir_data_in_1_), 
	.A0(FE_OFN517_n4693));
   AO22XLTS U2213 (.Y(n6363), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[4] ), 
	.B0(FE_OFN445_n4694), 
	.A1(FE_OFN1785_acc_fir_data_in_4_), 
	.A0(FE_OFN516_n4693));
   AO22XLTS U2208 (.Y(n6358), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[9] ), 
	.B0(FE_OFN446_n4694), 
	.A1(FE_OFN1755_acc_fir_data_in_9_), 
	.A0(FE_OFN520_n4693));
   AO22XLTS U2202 (.Y(n6352), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[15] ), 
	.B0(FE_OFN447_n4694), 
	.A1(FE_OFN1720_acc_fir_data_in_15_), 
	.A0(FE_OFN521_n4693));
   AO22XLTS U2210 (.Y(n6360), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[7] ), 
	.B0(FE_OFN448_n4694), 
	.A1(FE_OFN1768_acc_fir_data_in_7_), 
	.A0(FE_OFN515_n4693));
   AO22XLTS U1568 (.Y(n5820), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[18] ), 
	.B0(FE_OFN108_n4508), 
	.A1(FE_OFN1525_acc_fft_data_in_18_), 
	.A0(FE_OFN181_n4507));
   AO22XLTS U2191 (.Y(n6341), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[26] ), 
	.B0(FE_OFN451_n4694), 
	.A1(FE_OFN1657_acc_fir_data_in_26_), 
	.A0(FE_OFN512_n4693));
   AO22XLTS U2190 (.Y(n6340), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[27] ), 
	.B0(FE_OFN450_n4694), 
	.A1(FE_OFN1653_acc_fir_data_in_27_), 
	.A0(FE_OFN513_n4693));
   AO22XLTS U2212 (.Y(n6362), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[5] ), 
	.B0(FE_OFN450_n4694), 
	.A1(FE_OFN1782_acc_fir_data_in_5_), 
	.A0(FE_OFN515_n4693));
   AO22XLTS U2215 (.Y(n6365), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[2] ), 
	.B0(FE_OFN448_n4694), 
	.A1(FE_OFN1801_acc_fir_data_in_2_), 
	.A0(FE_OFN515_n4693));
   AO22XLTS U2204 (.Y(n6354), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[13] ), 
	.B0(FE_OFN446_n4694), 
	.A1(FE_OFN1735_acc_fir_data_in_13_), 
	.A0(FE_OFN520_n4693));
   AO22XLTS U2193 (.Y(n6343), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[24] ), 
	.B0(FE_OFN451_n4694), 
	.A1(FE_OFN1670_acc_fir_data_in_24_), 
	.A0(FE_OFN512_n4693));
   AO22XLTS U2192 (.Y(n6342), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[25] ), 
	.B0(FE_OFN451_n4694), 
	.A1(FE_OFN1665_acc_fir_data_in_25_), 
	.A0(FE_OFN512_n4693));
   AO22XLTS U1570 (.Y(n5822), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[16] ), 
	.B0(FE_OFN110_n4508), 
	.A1(FE_OFN1537_acc_fft_data_in_16_), 
	.A0(FE_OFN180_n4507));
   AO22XLTS U2207 (.Y(n6357), 
	.B1(\fifo_from_fir/fifo_cell12/sr_out[10] ), 
	.B0(FE_OFN447_n4694), 
	.A1(FE_OFN1747_acc_fir_data_in_10_), 
	.A0(FE_OFN521_n4693));
   AO22XLTS U1583 (.Y(n5835), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[3] ), 
	.B0(FE_OFN109_n4508), 
	.A1(FE_OFN1605_acc_fft_data_in_3_), 
	.A0(FE_OFN182_n4507));
   AO22XLTS U1585 (.Y(n5837), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[1] ), 
	.B0(FE_OFN107_n4508), 
	.A1(FE_OFN1617_acc_fft_data_in_1_), 
	.A0(FE_OFN179_n4507));
   AO22XLTS U1582 (.Y(n5834), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[4] ), 
	.B0(n4508), 
	.A1(FE_OFN1601_acc_fft_data_in_4_), 
	.A0(FE_OFN176_n4507));
   AO22XLTS U1586 (.Y(n5838), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[0] ), 
	.B0(FE_OFN109_n4508), 
	.A1(FE_OFN1624_acc_fft_data_in_0_), 
	.A0(FE_OFN182_n4507));
   AO22XLTS U1576 (.Y(n5828), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[10] ), 
	.B0(FE_OFN114_n4508), 
	.A1(FE_OFN1568_acc_fft_data_in_10_), 
	.A0(FE_OFN186_n4507));
   AO22XLTS U1575 (.Y(n5827), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[11] ), 
	.B0(FE_OFN114_n4508), 
	.A1(FE_OFN1559_acc_fft_data_in_11_), 
	.A0(FE_OFN186_n4507));
   AO22XLTS U1560 (.Y(n5812), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[26] ), 
	.B0(FE_OFN109_n4508), 
	.A1(FE_OFN1480_acc_fft_data_in_26_), 
	.A0(FE_OFN179_n4507));
   AO22XLTS U1577 (.Y(n5829), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[9] ), 
	.B0(FE_OFN114_n4508), 
	.A1(FE_OFN1571_acc_fft_data_in_9_), 
	.A0(FE_OFN186_n4507));
   AO22XLTS U1580 (.Y(n5832), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[6] ), 
	.B0(FE_OFN106_n4508), 
	.A1(FE_OFN1590_acc_fft_data_in_6_), 
	.A0(FE_OFN177_n4507));
   OAI21XLTS U2184 (.Y(n4689), 
	.B0(n8376), 
	.A1(n4692), 
	.A0(n7539));
   AO22XLTS U1574 (.Y(n5826), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[12] ), 
	.B0(FE_OFN112_n4508), 
	.A1(FE_OFN1553_acc_fft_data_in_12_), 
	.A0(FE_OFN183_n4507));
   AO22XLTS U1559 (.Y(n5811), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[27] ), 
	.B0(FE_OFN107_n4508), 
	.A1(FE_OFN1475_acc_fft_data_in_27_), 
	.A0(FE_OFN179_n4507));
   AO22XLTS U1573 (.Y(n5825), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[13] ), 
	.B0(FE_OFN110_n4508), 
	.A1(FE_OFN1548_acc_fft_data_in_13_), 
	.A0(FE_OFN181_n4507));
   AO22XLTS U1561 (.Y(n5813), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[25] ), 
	.B0(FE_OFN105_n4508), 
	.A1(FE_OFN1486_acc_fft_data_in_25_), 
	.A0(FE_OFN178_n4507));
   AO22XLTS U1579 (.Y(n5831), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[7] ), 
	.B0(FE_OFN106_n4508), 
	.A1(FE_OFN1582_acc_fft_data_in_7_), 
	.A0(FE_OFN177_n4507));
   AO22XLTS U1584 (.Y(n5836), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[2] ), 
	.B0(FE_OFN107_n4508), 
	.A1(FE_OFN1610_acc_fft_data_in_2_), 
	.A0(FE_OFN178_n4507));
   AO22XLTS U1572 (.Y(n5824), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[14] ), 
	.B0(FE_OFN112_n4508), 
	.A1(FE_OFN1543_acc_fft_data_in_14_), 
	.A0(FE_OFN183_n4507));
   AO22XLTS U1562 (.Y(n5814), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[24] ), 
	.B0(FE_OFN105_n4508), 
	.A1(FE_OFN1489_acc_fft_data_in_24_), 
	.A0(FE_OFN178_n4507));
   AO22XLTS U1581 (.Y(n5833), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[5] ), 
	.B0(FE_OFN106_n4508), 
	.A1(FE_OFN1595_acc_fft_data_in_5_), 
	.A0(FE_OFN177_n4507));
   AO22XLTS U1571 (.Y(n5823), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[15] ), 
	.B0(FE_OFN112_n4508), 
	.A1(FE_OFN1538_acc_fft_data_in_15_), 
	.A0(FE_OFN183_n4507));
   AO22XLTS U1578 (.Y(n5830), 
	.B1(\fifo_from_fft/fifo_cell12/sr_out[8] ), 
	.B0(FE_OFN114_n4508), 
	.A1(FE_OFN1579_acc_fft_data_in_8_), 
	.A0(FE_OFN186_n4507));
   NAND3XLTS U2658 (.Y(n4669), 
	.C(n4790), 
	.B(n4670), 
	.A(n8376));
   AO22XLTS U2158 (.Y(n6311), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[22] ), 
	.B0(FE_OFN462_n4688), 
	.A1(FE_OFN1679_acc_fir_data_in_22_), 
	.A0(n8382));
   OAI21XLTS U2183 (.Y(n6335), 
	.B0(n4689), 
	.A1(n4691), 
	.A0(\fifo_from_fir/fifo_cell13/data_out/N35 ));
   OAI21XLTS U1553 (.Y(n4503), 
	.B0(n8711), 
	.A1(n4506), 
	.A0(n7465));
   AO22XLTS U2159 (.Y(n6312), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[21] ), 
	.B0(FE_OFN462_n4688), 
	.A1(FE_OFN1685_acc_fir_data_in_21_), 
	.A0(n8382));
   AO22XLTS U2157 (.Y(n6310), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[23] ), 
	.B0(FE_OFN462_n4688), 
	.A1(FE_OFN1677_acc_fir_data_in_23_), 
	.A0(n8382));
   AO22XLTS U1527 (.Y(n5782), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[22] ), 
	.B0(FE_OFN123_n4502), 
	.A1(FE_OFN1504_acc_fft_data_in_22_), 
	.A0(n8717));
   AO22XLTS U2151 (.Y(n6304), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[29] ), 
	.B0(FE_OFN455_n4688), 
	.A1(FE_OFN1644_acc_fir_data_in_29_), 
	.A0(n8384));
   NAND3XLTS U2027 (.Y(n4483), 
	.C(n4604), 
	.B(n4484), 
	.A(n8711));
   AO22XLTS U2162 (.Y(n6315), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[18] ), 
	.B0(FE_OFN459_n4688), 
	.A1(FE_OFN1706_acc_fir_data_in_18_), 
	.A0(n8381));
   AO22XLTS U2163 (.Y(n6316), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[17] ), 
	.B0(FE_OFN458_n4688), 
	.A1(FE_OFN1711_acc_fir_data_in_17_), 
	.A0(n8381));
   AO22XLTS U2150 (.Y(n6303), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[30] ), 
	.B0(FE_OFN455_n4688), 
	.A1(FE_OFN1636_acc_fir_data_in_30_), 
	.A0(n8384));
   AO22XLTS U2161 (.Y(n6314), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[19] ), 
	.B0(FE_OFN458_n4688), 
	.A1(FE_OFN1697_acc_fir_data_in_19_), 
	.A0(n8381));
   AO22XLTS U2164 (.Y(n6317), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[16] ), 
	.B0(FE_OFN458_n4688), 
	.A1(FE_OFN1718_acc_fir_data_in_16_), 
	.A0(n8381));
   OAI211XLTS U2659 (.Y(n4789), 
	.C0(n9468), 
	.B0(\fifo_from_fir/hang[12] ), 
	.A1(n4791), 
	.A0(n8874));
   OAI21XLTS U1552 (.Y(n5806), 
	.B0(n4503), 
	.A1(n4505), 
	.A0(\fifo_from_fft/fifo_cell13/data_out/N35 ));
   AO22XLTS U2149 (.Y(n6302), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[31] ), 
	.B0(FE_OFN455_n4688), 
	.A1(FE_OFN1631_acc_fir_data_in_31_), 
	.A0(n8384));
   AO22XLTS U2160 (.Y(n6313), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[20] ), 
	.B0(FE_OFN462_n4688), 
	.A1(FE_OFN1694_acc_fir_data_in_20_), 
	.A0(n8382));
   AO22XLTS U2152 (.Y(n6305), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[28] ), 
	.B0(FE_OFN455_n4688), 
	.A1(FE_OFN1649_acc_fir_data_in_28_), 
	.A0(n8384));
   AO22XLTS U1518 (.Y(n5773), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[31] ), 
	.B0(FE_OFN118_n4502), 
	.A1(FE_OFN1456_acc_fft_data_in_31_), 
	.A0(n8719));
   OAI211XLTS U2028 (.Y(n4603), 
	.C0(n9470), 
	.B0(\fifo_from_fft/hang[12] ), 
	.A1(n4605), 
	.A0(n8841));
   AO22XLTS U1526 (.Y(n5781), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[23] ), 
	.B0(FE_OFN124_n4502), 
	.A1(FE_OFN1495_acc_fft_data_in_23_), 
	.A0(n8717));
   AO22XLTS U1531 (.Y(n5786), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[18] ), 
	.B0(FE_OFN128_n4502), 
	.A1(FE_OFN1526_acc_fft_data_in_18_), 
	.A0(n8716));
   AO22XLTS U1530 (.Y(n5785), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[19] ), 
	.B0(FE_OFN128_n4502), 
	.A1(FE_OFN1515_acc_fft_data_in_19_), 
	.A0(n8716));
   AO22XLTS U1533 (.Y(n5788), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[16] ), 
	.B0(FE_OFN128_n4502), 
	.A1(FE_OFN1535_acc_fft_data_in_16_), 
	.A0(n8716));
   AO22XLTS U1519 (.Y(n5774), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[30] ), 
	.B0(FE_OFN118_n4502), 
	.A1(FE_OFN1462_acc_fft_data_in_30_), 
	.A0(n8719));
   AO22XLTS U1520 (.Y(n5775), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[29] ), 
	.B0(FE_OFN118_n4502), 
	.A1(FE_OFN1467_acc_fft_data_in_29_), 
	.A0(n8719));
   AO22XLTS U1532 (.Y(n5787), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[17] ), 
	.B0(FE_OFN128_n4502), 
	.A1(FE_OFN1532_acc_fft_data_in_17_), 
	.A0(n8716));
   AO22XLTS U1529 (.Y(n5784), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[20] ), 
	.B0(FE_OFN124_n4502), 
	.A1(FE_OFN1513_acc_fft_data_in_20_), 
	.A0(n8717));
   AO22XLTS U1528 (.Y(n5783), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[21] ), 
	.B0(FE_OFN123_n4502), 
	.A1(FE_OFN1508_acc_fft_data_in_21_), 
	.A0(n8717));
   AO22XLTS U2153 (.Y(n6306), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[27] ), 
	.B0(FE_OFN453_n4688), 
	.A1(FE_OFN1654_acc_fir_data_in_27_), 
	.A0(n8383));
   AO22XLTS U2156 (.Y(n6309), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[24] ), 
	.B0(FE_OFN453_n4688), 
	.A1(FE_OFN1668_acc_fir_data_in_24_), 
	.A0(n8383));
   AO22XLTS U2174 (.Y(n6327), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[6] ), 
	.B0(FE_OFN454_n4688), 
	.A1(FE_OFN1776_acc_fir_data_in_6_), 
	.A0(n8378));
   AO22XLTS U2179 (.Y(n6332), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[1] ), 
	.B0(FE_OFN457_n4688), 
	.A1(FE_OFN1802_acc_fir_data_in_1_), 
	.A0(n8377));
   AO22XLTS U2173 (.Y(n6326), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[7] ), 
	.B0(FE_OFN454_n4688), 
	.A1(FE_OFN1768_acc_fir_data_in_7_), 
	.A0(n8378));
   AO22XLTS U2176 (.Y(n6329), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[4] ), 
	.B0(FE_OFN454_n4688), 
	.A1(FE_OFN1789_acc_fir_data_in_4_), 
	.A0(n8378));
   AO22XLTS U2154 (.Y(n6307), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[26] ), 
	.B0(FE_OFN453_n4688), 
	.A1(FE_OFN1660_acc_fir_data_in_26_), 
	.A0(n8383));
   AO22XLTS U2168 (.Y(n6321), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[12] ), 
	.B0(FE_OFN460_n4688), 
	.A1(FE_OFN1740_acc_fir_data_in_12_), 
	.A0(n8380));
   AO22XLTS U2167 (.Y(n6320), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[13] ), 
	.B0(FE_OFN459_n4688), 
	.A1(FE_OFN1735_acc_fir_data_in_13_), 
	.A0(n8380));
   AO22XLTS U2172 (.Y(n6325), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[8] ), 
	.B0(FE_OFN461_n4688), 
	.A1(FE_OFN1758_acc_fir_data_in_8_), 
	.A0(n8379));
   AO22XLTS U2177 (.Y(n6330), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[3] ), 
	.B0(FE_OFN457_n4688), 
	.A1(FE_OFN1792_acc_fir_data_in_3_), 
	.A0(n8377));
   AO22XLTS U2155 (.Y(n6308), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[25] ), 
	.B0(n4688), 
	.A1(FE_OFN1662_acc_fir_data_in_25_), 
	.A0(n8383));
   AO22XLTS U2169 (.Y(n6322), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[11] ), 
	.B0(FE_OFN461_n4688), 
	.A1(FE_OFN1743_acc_fir_data_in_11_), 
	.A0(n8379));
   AO22XLTS U2180 (.Y(n6333), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[0] ), 
	.B0(FE_OFN457_n4688), 
	.A1(FE_OFN1814_acc_fir_data_in_0_), 
	.A0(n8377));
   AO22XLTS U2178 (.Y(n6331), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[2] ), 
	.B0(FE_OFN456_n4688), 
	.A1(FE_OFN1799_acc_fir_data_in_2_), 
	.A0(n8377));
   AO22XLTS U2175 (.Y(n6328), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[5] ), 
	.B0(n4688), 
	.A1(FE_OFN1779_acc_fir_data_in_5_), 
	.A0(n8378));
   AO22XLTS U2165 (.Y(n6318), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[15] ), 
	.B0(FE_OFN460_n4688), 
	.A1(FE_OFN1722_acc_fir_data_in_15_), 
	.A0(n8380));
   AO22XLTS U2171 (.Y(n6324), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[9] ), 
	.B0(FE_OFN461_n4688), 
	.A1(FE_OFN1755_acc_fir_data_in_9_), 
	.A0(n8379));
   AO22XLTS U1521 (.Y(n5776), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[28] ), 
	.B0(FE_OFN116_n4502), 
	.A1(FE_OFN1471_acc_fft_data_in_28_), 
	.A0(n8719));
   AO22XLTS U2166 (.Y(n6319), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[14] ), 
	.B0(FE_OFN460_n4688), 
	.A1(FE_OFN1729_acc_fir_data_in_14_), 
	.A0(n8380));
   AO22XLTS U2170 (.Y(n6323), 
	.B1(\fifo_from_fir/fifo_cell13/sr_out[10] ), 
	.B0(FE_OFN461_n4688), 
	.A1(FE_OFN1750_acc_fir_data_in_10_), 
	.A0(n8379));
   AO22XLTS U1538 (.Y(n5793), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[11] ), 
	.B0(FE_OFN125_n4502), 
	.A1(FE_OFN1562_acc_fft_data_in_11_), 
	.A0(n8714));
   AO22XLTS U1522 (.Y(n5777), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[27] ), 
	.B0(FE_OFN122_n4502), 
	.A1(FE_OFN1477_acc_fft_data_in_27_), 
	.A0(n8718));
   AO22XLTS U1523 (.Y(n5778), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[26] ), 
	.B0(FE_OFN122_n4502), 
	.A1(FE_OFN1482_acc_fft_data_in_26_), 
	.A0(n8718));
   AO22XLTS U1524 (.Y(n5779), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[25] ), 
	.B0(FE_OFN120_n4502), 
	.A1(FE_OFN1487_acc_fft_data_in_25_), 
	.A0(n8718));
   AO22XLTS U1545 (.Y(n5800), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[4] ), 
	.B0(n4502), 
	.A1(FE_OFN1602_acc_fft_data_in_4_), 
	.A0(n8713));
   AO22XLTS U1544 (.Y(n5799), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[5] ), 
	.B0(FE_OFN116_n4502), 
	.A1(FE_OFN1595_acc_fft_data_in_5_), 
	.A0(n8713));
   AO22XLTS U1542 (.Y(n5797), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[7] ), 
	.B0(FE_OFN115_n4502), 
	.A1(FE_OFN1580_acc_fft_data_in_7_), 
	.A0(n8713));
   AO22XLTS U1543 (.Y(n5798), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[6] ), 
	.B0(FE_OFN115_n4502), 
	.A1(FE_OFN1590_acc_fft_data_in_6_), 
	.A0(n8713));
   AO22XLTS U1540 (.Y(n5795), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[9] ), 
	.B0(FE_OFN125_n4502), 
	.A1(FE_OFN1572_acc_fft_data_in_9_), 
	.A0(n8714));
   AO22XLTS U1537 (.Y(n5792), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[12] ), 
	.B0(FE_OFN127_n4502), 
	.A1(FE_OFN1557_acc_fft_data_in_12_), 
	.A0(n8715));
   AO22XLTS U1547 (.Y(n5802), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[2] ), 
	.B0(FE_OFN119_n4502), 
	.A1(FE_OFN1613_acc_fft_data_in_2_), 
	.A0(n8712));
   AO22XLTS U1536 (.Y(n5791), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[13] ), 
	.B0(FE_OFN126_n4502), 
	.A1(FE_OFN1552_acc_fft_data_in_13_), 
	.A0(n8715));
   AO22XLTS U1535 (.Y(n5790), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[14] ), 
	.B0(FE_OFN127_n4502), 
	.A1(FE_OFN1545_acc_fft_data_in_14_), 
	.A0(n8715));
   AO22XLTS U1539 (.Y(n5794), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[10] ), 
	.B0(FE_OFN125_n4502), 
	.A1(FE_OFN1567_acc_fft_data_in_10_), 
	.A0(n8714));
   AO22XLTS U1549 (.Y(n5804), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[0] ), 
	.B0(FE_OFN122_n4502), 
	.A1(FE_OFN1626_acc_fft_data_in_0_), 
	.A0(n8712));
   AO22XLTS U1534 (.Y(n5789), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[15] ), 
	.B0(FE_OFN126_n4502), 
	.A1(FE_OFN1541_acc_fft_data_in_15_), 
	.A0(n8715));
   AO22XLTS U1546 (.Y(n5801), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[3] ), 
	.B0(FE_OFN122_n4502), 
	.A1(FE_OFN1606_acc_fft_data_in_3_), 
	.A0(n8712));
   AO22XLTS U1541 (.Y(n5796), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[8] ), 
	.B0(FE_OFN126_n4502), 
	.A1(FE_OFN1576_acc_fft_data_in_8_), 
	.A0(n8714));
   AO22XLTS U1525 (.Y(n5780), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[24] ), 
	.B0(FE_OFN120_n4502), 
	.A1(FE_OFN1492_acc_fft_data_in_24_), 
	.A0(n8718));
   AO22XLTS U1548 (.Y(n5803), 
	.B1(\fifo_from_fft/fifo_cell13/sr_out[1] ), 
	.B0(FE_OFN119_n4502), 
	.A1(FE_OFN1621_acc_fft_data_in_1_), 
	.A0(n8712));
   OAI21XLTS U2147 (.Y(n4683), 
	.B0(FE_OFN496_n4681), 
	.A1(n4686), 
	.A0(n7534));
   OAI21X1TS U1516 (.Y(n4497), 
	.B0(FE_OFN161_n4495), 
	.A1(n4500), 
	.A0(n7460));
   OAI21XLTS U2146 (.Y(n6301), 
	.B0(n4683), 
	.A1(n4685), 
	.A0(\fifo_from_fir/fifo_cell14/data_out/N35 ));
   NAND3XLTS U2656 (.Y(n4671), 
	.C(n4787), 
	.B(n4672), 
	.A(FE_OFN496_n4681));
   AO22XLTS U2122 (.Y(n6278), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[21] ), 
	.B0(FE_OFN486_n4682), 
	.A1(FE_OFN1689_acc_fir_data_in_21_), 
	.A0(FE_OFN504_n4681));
   OAI211XLTS U2657 (.Y(n4786), 
	.C0(n9469), 
	.B0(\fifo_from_fir/hang[13] ), 
	.A1(n4788), 
	.A0(n8874));
   AO22XLTS U2138 (.Y(n6294), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[5] ), 
	.B0(FE_OFN490_n4682), 
	.A1(FE_OFN1778_acc_fir_data_in_5_), 
	.A0(FE_OFN500_n4681));
   OAI21XLTS U1515 (.Y(n5772), 
	.B0(n4497), 
	.A1(n4499), 
	.A0(\fifo_from_fft/fifo_cell14/data_out/N35 ));
   AO22XLTS U2137 (.Y(n6293), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[6] ), 
	.B0(FE_OFN492_n4682), 
	.A1(FE_OFN1775_acc_fir_data_in_6_), 
	.A0(FE_OFN500_n4681));
   AO22XLTS U2136 (.Y(n6292), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[7] ), 
	.B0(FE_OFN490_n4682), 
	.A1(FE_OFN1762_acc_fir_data_in_7_), 
	.A0(FE_OFN500_n4681));
   AO22XLTS U2139 (.Y(n6295), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[4] ), 
	.B0(FE_OFN488_n4682), 
	.A1(FE_OFN1788_acc_fir_data_in_4_), 
	.A0(FE_OFN501_n4681));
   NAND3XLTS U2025 (.Y(n4485), 
	.C(n4601), 
	.B(n4486), 
	.A(n4495));
   AO22XLTS U1491 (.Y(n5749), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[21] ), 
	.B0(FE_OFN157_n4496), 
	.A1(FE_OFN1507_acc_fft_data_in_21_), 
	.A0(FE_OFN171_n4495));
   AO22XLTS U2112 (.Y(n6268), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[31] ), 
	.B0(FE_OFN493_n4682), 
	.A1(FE_OFN1628_acc_fir_data_in_31_), 
	.A0(FE_OFN499_n4681));
   AO22XLTS U2113 (.Y(n6269), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[30] ), 
	.B0(FE_OFN492_n4682), 
	.A1(FE_OFN1635_acc_fir_data_in_30_), 
	.A0(FE_OFN498_n4681));
   AO22XLTS U2120 (.Y(n6276), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[23] ), 
	.B0(FE_OFN487_n4682), 
	.A1(FE_OFN1671_acc_fir_data_in_23_), 
	.A0(FE_OFN503_n4681));
   AO22XLTS U2121 (.Y(n6277), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[22] ), 
	.B0(FE_OFN486_n4682), 
	.A1(FE_OFN1679_acc_fir_data_in_22_), 
	.A0(FE_OFN504_n4681));
   AO22XLTS U2123 (.Y(n6279), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[20] ), 
	.B0(FE_OFN487_n4682), 
	.A1(FE_OFN1691_acc_fir_data_in_20_), 
	.A0(FE_OFN504_n4681));
   AO22XLTS U2114 (.Y(n6270), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[29] ), 
	.B0(FE_OFN493_n4682), 
	.A1(FE_OFN1638_acc_fir_data_in_29_), 
	.A0(FE_OFN499_n4681));
   AO22XLTS U1481 (.Y(n5739), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[31] ), 
	.B0(FE_OFN157_n4496), 
	.A1(FE_OFN1453_acc_fft_data_in_31_), 
	.A0(FE_OFN171_n4495));
   OAI211XLTS U2026 (.Y(n4600), 
	.C0(n9472), 
	.B0(\fifo_from_fft/hang[13] ), 
	.A1(n4602), 
	.A0(n8841));
   AO22XLTS U1482 (.Y(n5740), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[30] ), 
	.B0(FE_OFN155_n4496), 
	.A1(FE_OFN1460_acc_fft_data_in_30_), 
	.A0(FE_OFN170_n4495));
   AO22XLTS U1490 (.Y(n5748), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[22] ), 
	.B0(FE_OFN157_n4496), 
	.A1(FE_OFN1501_acc_fft_data_in_22_), 
	.A0(FE_OFN171_n4495));
   AO22XLTS U1489 (.Y(n5747), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[23] ), 
	.B0(FE_OFN154_n4496), 
	.A1(FE_OFN1495_acc_fft_data_in_23_), 
	.A0(FE_OFN169_n4495));
   AO22XLTS U1483 (.Y(n5741), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[29] ), 
	.B0(FE_OFN155_n4496), 
	.A1(FE_OFN1466_acc_fft_data_in_29_), 
	.A0(FE_OFN170_n4495));
   AO22XLTS U1492 (.Y(n5750), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[20] ), 
	.B0(FE_OFN154_n4496), 
	.A1(FE_OFN1512_acc_fft_data_in_20_), 
	.A0(FE_OFN169_n4495));
   AO22XLTS U1507 (.Y(n5765), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[5] ), 
	.B0(FE_OFN154_n4496), 
	.A1(FE_OFN1592_acc_fft_data_in_5_), 
	.A0(FE_OFN166_n4495));
   AO22XLTS U1506 (.Y(n5764), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[6] ), 
	.B0(FE_OFN156_n4496), 
	.A1(FE_OFN1589_acc_fft_data_in_6_), 
	.A0(FE_OFN169_n4495));
   AO22XLTS U1505 (.Y(n5763), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[7] ), 
	.B0(FE_OFN151_n4496), 
	.A1(FE_OFN1583_acc_fft_data_in_7_), 
	.A0(FE_OFN164_n4495));
   AO22XLTS U1508 (.Y(n5766), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[4] ), 
	.B0(FE_OFN158_n4496), 
	.A1(FE_OFN1599_acc_fft_data_in_4_), 
	.A0(FE_OFN163_n4495));
   AO22XLTS U2115 (.Y(n6271), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[28] ), 
	.B0(FE_OFN493_n4682), 
	.A1(FE_OFN1646_acc_fir_data_in_28_), 
	.A0(FE_OFN499_n4681));
   AO22XLTS U2141 (.Y(n6297), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[2] ), 
	.B0(FE_OFN488_n4682), 
	.A1(FE_OFN1796_acc_fir_data_in_2_), 
	.A0(FE_OFN501_n4681));
   AO22XLTS U2124 (.Y(n6280), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[19] ), 
	.B0(FE_OFN487_n4682), 
	.A1(FE_OFN1698_acc_fir_data_in_19_), 
	.A0(FE_OFN503_n4681));
   AO22XLTS U2142 (.Y(n6298), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[1] ), 
	.B0(n4682), 
	.A1(FE_OFN1805_acc_fir_data_in_1_), 
	.A0(FE_OFN502_n4681));
   AO22XLTS U2135 (.Y(n6291), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[8] ), 
	.B0(FE_OFN495_n4682), 
	.A1(FE_OFN1757_acc_fir_data_in_8_), 
	.A0(FE_OFN507_n4681));
   AO22XLTS U2126 (.Y(n6282), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[17] ), 
	.B0(FE_OFN491_n4682), 
	.A1(FE_OFN1710_acc_fir_data_in_17_), 
	.A0(FE_OFN505_n4681));
   AO22XLTS U2125 (.Y(n6281), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[18] ), 
	.B0(FE_OFN491_n4682), 
	.A1(FE_OFN1702_acc_fir_data_in_18_), 
	.A0(FE_OFN505_n4681));
   AO22XLTS U2117 (.Y(n6273), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[26] ), 
	.B0(FE_OFN494_n4682), 
	.A1(FE_OFN1658_acc_fir_data_in_26_), 
	.A0(FE_OFN498_n4681));
   AO22XLTS U2127 (.Y(n6283), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[16] ), 
	.B0(FE_OFN491_n4682), 
	.A1(FE_OFN1712_acc_fir_data_in_16_), 
	.A0(FE_OFN505_n4681));
   AO22XLTS U2116 (.Y(n6272), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[27] ), 
	.B0(FE_OFN494_n4682), 
	.A1(FE_OFN1651_acc_fir_data_in_27_), 
	.A0(FE_OFN498_n4681));
   AO22XLTS U2140 (.Y(n6296), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[3] ), 
	.B0(n4682), 
	.A1(FE_OFN1794_acc_fir_data_in_3_), 
	.A0(FE_OFN502_n4681));
   AO22XLTS U2128 (.Y(n6284), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[15] ), 
	.B0(FE_OFN489_n4682), 
	.A1(FE_OFN1722_acc_fir_data_in_15_), 
	.A0(FE_OFN506_n4681));
   AO22XLTS U2129 (.Y(n6285), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[14] ), 
	.B0(FE_OFN489_n4682), 
	.A1(FE_OFN1729_acc_fir_data_in_14_), 
	.A0(FE_OFN506_n4681));
   AO22XLTS U2132 (.Y(n6288), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[11] ), 
	.B0(FE_OFN495_n4682), 
	.A1(FE_OFN1741_acc_fir_data_in_11_), 
	.A0(FE_OFN507_n4681));
   AO22XLTS U2143 (.Y(n6299), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[0] ), 
	.B0(FE_OFN488_n4682), 
	.A1(FE_OFN1812_acc_fir_data_in_0_), 
	.A0(FE_OFN501_n4681));
   AO22XLTS U1484 (.Y(n5742), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[28] ), 
	.B0(FE_OFN155_n4496), 
	.A1(FE_OFN1470_acc_fft_data_in_28_), 
	.A0(FE_OFN170_n4495));
   AO22XLTS U2118 (.Y(n6274), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[25] ), 
	.B0(FE_OFN494_n4682), 
	.A1(FE_OFN1664_acc_fir_data_in_25_), 
	.A0(FE_OFN497_n4681));
   AO22XLTS U2133 (.Y(n6289), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[10] ), 
	.B0(FE_OFN489_n4682), 
	.A1(FE_OFN1750_acc_fir_data_in_10_), 
	.A0(FE_OFN506_n4681));
   AO22XLTS U2134 (.Y(n6290), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[9] ), 
	.B0(FE_OFN495_n4682), 
	.A1(FE_OFN1753_acc_fir_data_in_9_), 
	.A0(FE_OFN507_n4681));
   AO22XLTS U2119 (.Y(n6275), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[24] ), 
	.B0(FE_OFN494_n4682), 
	.A1(FE_OFN1669_acc_fir_data_in_24_), 
	.A0(FE_OFN497_n4681));
   AO22XLTS U2131 (.Y(n6287), 
	.B1(\fifo_from_fir/fifo_cell14/sr_out[12] ), 
	.B0(FE_OFN489_n4682), 
	.A1(FE_OFN1740_acc_fir_data_in_12_), 
	.A0(FE_OFN506_n4681));
   AO22XLTS U1503 (.Y(n5761), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[9] ), 
	.B0(FE_OFN160_n4496), 
	.A1(FE_OFN1573_acc_fft_data_in_9_), 
	.A0(FE_OFN172_n4495));
   AO22XLTS U1495 (.Y(n5753), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[17] ), 
	.B0(FE_OFN158_n4496), 
	.A1(FE_OFN1530_acc_fft_data_in_17_), 
	.A0(FE_OFN165_n4495));
   AO22XLTS U1496 (.Y(n5754), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[16] ), 
	.B0(FE_OFN158_n4496), 
	.A1(FE_OFN1535_acc_fft_data_in_16_), 
	.A0(FE_OFN165_n4495));
   AO22XLTS U1501 (.Y(n5759), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[11] ), 
	.B0(FE_OFN160_n4496), 
	.A1(FE_OFN1560_acc_fft_data_in_11_), 
	.A0(FE_OFN172_n4495));
   AO22XLTS U1494 (.Y(n5752), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[18] ), 
	.B0(FE_OFN156_n4496), 
	.A1(FE_OFN1525_acc_fft_data_in_18_), 
	.A0(FE_OFN169_n4495));
   AO22XLTS U1497 (.Y(n5755), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[15] ), 
	.B0(FE_OFN159_n4496), 
	.A1(FE_OFN1539_acc_fft_data_in_15_), 
	.A0(FE_OFN167_n4495));
   AO22XLTS U1498 (.Y(n5756), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[14] ), 
	.B0(FE_OFN159_n4496), 
	.A1(FE_OFN1545_acc_fft_data_in_14_), 
	.A0(FE_OFN167_n4495));
   AO22XLTS U1493 (.Y(n5751), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[19] ), 
	.B0(FE_OFN158_n4496), 
	.A1(FE_OFN1517_acc_fft_data_in_19_), 
	.A0(FE_OFN163_n4495));
   AO22XLTS U1502 (.Y(n5760), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[10] ), 
	.B0(FE_OFN160_n4496), 
	.A1(FE_OFN1565_acc_fft_data_in_10_), 
	.A0(FE_OFN172_n4495));
   AO22XLTS U1500 (.Y(n5758), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[12] ), 
	.B0(FE_OFN159_n4496), 
	.A1(FE_OFN1554_acc_fft_data_in_12_), 
	.A0(FE_OFN165_n4495));
   AO22XLTS U1504 (.Y(n5762), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[8] ), 
	.B0(FE_OFN160_n4496), 
	.A1(FE_OFN1578_acc_fft_data_in_8_), 
	.A0(FE_OFN172_n4495));
   AO22XLTS U1487 (.Y(n5745), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[25] ), 
	.B0(n4496), 
	.A1(FE_OFN1484_acc_fft_data_in_25_), 
	.A0(FE_OFN162_n4495));
   AO22XLTS U1510 (.Y(n5768), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[2] ), 
	.B0(FE_OFN151_n4496), 
	.A1(FE_OFN1610_acc_fft_data_in_2_), 
	.A0(FE_OFN164_n4495));
   AO22XLTS U1509 (.Y(n5767), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[3] ), 
	.B0(FE_OFN153_n4496), 
	.A1(FE_OFN1604_acc_fft_data_in_3_), 
	.A0(FE_OFN168_n4495));
   AO22XLTS U1511 (.Y(n5769), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[1] ), 
	.B0(FE_OFN151_n4496), 
	.A1(FE_OFN1616_acc_fft_data_in_1_), 
	.A0(FE_OFN164_n4495));
   AO22XLTS U1485 (.Y(n5743), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[27] ), 
	.B0(FE_OFN152_n4496), 
	.A1(FE_OFN1474_acc_fft_data_in_27_), 
	.A0(FE_OFN166_n4495));
   AO22XLTS U1486 (.Y(n5744), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[26] ), 
	.B0(FE_OFN152_n4496), 
	.A1(FE_OFN1478_acc_fft_data_in_26_), 
	.A0(FE_OFN166_n4495));
   AO22XLTS U1512 (.Y(n5770), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[0] ), 
	.B0(FE_OFN153_n4496), 
	.A1(FE_OFN1623_acc_fft_data_in_0_), 
	.A0(FE_OFN168_n4495));
   AO22XLTS U1488 (.Y(n5746), 
	.B1(\fifo_from_fft/fifo_cell14/sr_out[24] ), 
	.B0(n4496), 
	.A1(FE_OFN1490_acc_fft_data_in_24_), 
	.A0(FE_OFN162_n4495));
   OAI21X1TS U2110 (.Y(n4677), 
	.B0(n4675), 
	.A1(n4680), 
	.A0(n7529));
   AO22XLTS U2102 (.Y(n6261), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[4] ), 
	.B0(FE_OFN465_n4676), 
	.A1(FE_OFN1786_acc_fir_data_in_4_), 
	.A0(FE_OFN478_n4675));
   NAND3XLTS U2654 (.Y(n4673), 
	.C(n4784), 
	.B(n4674), 
	.A(FE_OFN474_n4675));
   INVXLTS U3612 (.Y(n4785), 
	.A(n4674));
   OAI21XLTS U2109 (.Y(n6267), 
	.B0(n4677), 
	.A1(n4679), 
	.A0(\fifo_from_fir/fifo_cell15/data_out/N35 ));
   OAI21XLTS U1479 (.Y(n4491), 
	.B0(n4489), 
	.A1(n4494), 
	.A0(n7455));
   NAND3XLTS U2023 (.Y(n4487), 
	.C(n4598), 
	.B(n4488), 
	.A(n4489));
   OAI21XLTS U1478 (.Y(n5738), 
	.B0(n4491), 
	.A1(n4493), 
	.A0(\fifo_from_fft/fifo_cell15/data_out/N35 ));
   INVXLTS U3755 (.Y(n4599), 
	.A(n4488));
   AO22XLTS U2101 (.Y(n6260), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[5] ), 
	.B0(FE_OFN467_n4676), 
	.A1(FE_OFN1781_acc_fir_data_in_5_), 
	.A0(FE_OFN475_n4675));
   AO22XLTS U1471 (.Y(n5732), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[4] ), 
	.B0(FE_OFN129_n4490), 
	.A1(FE_OFN1597_acc_fft_data_in_4_), 
	.A0(FE_OFN143_n4489));
   AO22XLTS U2100 (.Y(n6259), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[6] ), 
	.B0(FE_OFN465_n4676), 
	.A1(FE_OFN1770_acc_fir_data_in_6_), 
	.A0(FE_OFN478_n4675));
   AO22XLTS U2099 (.Y(n6258), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[7] ), 
	.B0(FE_OFN465_n4676), 
	.A1(FE_OFN1765_acc_fir_data_in_7_), 
	.A0(FE_OFN478_n4675));
   AO22XLTS U2096 (.Y(n6255), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[10] ), 
	.B0(FE_OFN471_n4676), 
	.A1(FE_OFN1746_acc_fir_data_in_10_), 
	.A0(FE_OFN483_n4675));
   AO22XLTS U2080 (.Y(n6239), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[26] ), 
	.B0(FE_OFN469_n4676), 
	.A1(FE_OFN1818_acc_fir_data_in_26_), 
	.A0(FE_OFN476_n4675));
   AO22XLTS U2097 (.Y(n6256), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[9] ), 
	.B0(FE_OFN472_n4676), 
	.A1(FE_OFN1755_acc_fir_data_in_9_), 
	.A0(FE_OFN484_n4675));
   AO22XLTS U2089 (.Y(n6248), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[17] ), 
	.B0(FE_OFN466_n4676), 
	.A1(FE_OFN1710_acc_fir_data_in_17_), 
	.A0(FE_OFN481_n4675));
   AO22XLTS U2076 (.Y(n6235), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[30] ), 
	.B0(FE_OFN470_n4676), 
	.A1(FE_OFN1633_acc_fir_data_in_30_), 
	.A0(FE_OFN476_n4675));
   AO22XLTS U2082 (.Y(n6241), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[24] ), 
	.B0(FE_OFN469_n4676), 
	.A1(FE_OFN1669_acc_fir_data_in_24_), 
	.A0(FE_OFN475_n4675));
   AO22XLTS U2075 (.Y(n6234), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[31] ), 
	.B0(FE_OFN470_n4676), 
	.A1(FE_OFN1632_acc_fir_data_in_31_), 
	.A0(FE_OFN477_n4675));
   AO22XLTS U2093 (.Y(n6252), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[13] ), 
	.B0(FE_OFN468_n4676), 
	.A1(FE_OFN1734_acc_fir_data_in_13_), 
	.A0(FE_OFN482_n4675));
   AO22XLTS U2084 (.Y(n6243), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[22] ), 
	.B0(FE_OFN473_n4676), 
	.A1(FE_OFN1680_acc_fir_data_in_22_), 
	.A0(FE_OFN485_n4675));
   AO22XLTS U2083 (.Y(n6242), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[23] ), 
	.B0(FE_OFN468_n4676), 
	.A1(FE_OFN1673_acc_fir_data_in_23_), 
	.A0(FE_OFN482_n4675));
   AO22XLTS U2086 (.Y(n6245), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[20] ), 
	.B0(n4676), 
	.A1(FE_OFN1693_acc_fir_data_in_20_), 
	.A0(FE_OFN480_n4675));
   AO22XLTS U1469 (.Y(n5730), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[6] ), 
	.B0(FE_OFN130_n4490), 
	.A1(FE_OFN1586_acc_fft_data_in_6_), 
	.A0(FE_OFN145_n4489));
   AO22XLTS U2094 (.Y(n6253), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[12] ), 
	.B0(FE_OFN473_n4676), 
	.A1(FE_OFN1737_acc_fir_data_in_12_), 
	.A0(FE_OFN485_n4675));
   AO22XLTS U2092 (.Y(n6251), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[14] ), 
	.B0(FE_OFN473_n4676), 
	.A1(FE_OFN1724_acc_fir_data_in_14_), 
	.A0(FE_OFN485_n4675));
   AO22XLTS U2085 (.Y(n6244), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[21] ), 
	.B0(FE_OFN473_n4676), 
	.A1(FE_OFN1688_acc_fir_data_in_21_), 
	.A0(FE_OFN485_n4675));
   AO22XLTS U2087 (.Y(n6246), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[19] ), 
	.B0(FE_OFN466_n4676), 
	.A1(FE_OFN1700_acc_fir_data_in_19_), 
	.A0(FE_OFN480_n4675));
   AO22XLTS U2081 (.Y(n6240), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[25] ), 
	.B0(FE_OFN469_n4676), 
	.A1(FE_OFN1664_acc_fir_data_in_25_), 
	.A0(FE_OFN475_n4675));
   AO22XLTS U1468 (.Y(n5729), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[7] ), 
	.B0(n4490), 
	.A1(FE_OFN1581_acc_fft_data_in_7_), 
	.A0(FE_OFN142_n4489));
   AO22XLTS U2103 (.Y(n6262), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[3] ), 
	.B0(FE_OFN464_n4676), 
	.A1(FE_OFN1791_acc_fir_data_in_3_), 
	.A0(FE_OFN479_n4675));
   AO22XLTS U2079 (.Y(n6238), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[27] ), 
	.B0(FE_OFN467_n4676), 
	.A1(FE_OFN1651_acc_fir_data_in_27_), 
	.A0(FE_OFN476_n4675));
   AO22XLTS U2091 (.Y(n6250), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[15] ), 
	.B0(FE_OFN471_n4676), 
	.A1(FE_OFN1719_acc_fir_data_in_15_), 
	.A0(FE_OFN483_n4675));
   AO22XLTS U2095 (.Y(n6254), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[11] ), 
	.B0(FE_OFN472_n4676), 
	.A1(FE_OFN1742_acc_fir_data_in_11_), 
	.A0(FE_OFN484_n4675));
   AO22XLTS U2088 (.Y(n6247), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[18] ), 
	.B0(FE_OFN468_n4676), 
	.A1(FE_OFN1705_acc_fir_data_in_18_), 
	.A0(FE_OFN482_n4675));
   AO22XLTS U2090 (.Y(n6249), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[16] ), 
	.B0(FE_OFN466_n4676), 
	.A1(FE_OFN1717_acc_fir_data_in_16_), 
	.A0(FE_OFN481_n4675));
   AO22XLTS U1470 (.Y(n5731), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[5] ), 
	.B0(FE_OFN131_n4490), 
	.A1(FE_OFN1591_acc_fft_data_in_5_), 
	.A0(FE_OFN145_n4489));
   AO22XLTS U2078 (.Y(n6237), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[28] ), 
	.B0(FE_OFN470_n4676), 
	.A1(FE_OFN1648_acc_fir_data_in_28_), 
	.A0(FE_OFN477_n4675));
   AO22XLTS U2106 (.Y(n6265), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[0] ), 
	.B0(FE_OFN464_n4676), 
	.A1(FE_OFN1808_acc_fir_data_in_0_), 
	.A0(FE_OFN481_n4675));
   AO22XLTS U2104 (.Y(n6263), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[2] ), 
	.B0(FE_OFN463_n4676), 
	.A1(FE_OFN1799_acc_fir_data_in_2_), 
	.A0(FE_OFN479_n4675));
   AO22XLTS U2098 (.Y(n6257), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[8] ), 
	.B0(FE_OFN472_n4676), 
	.A1(FE_OFN1760_acc_fir_data_in_8_), 
	.A0(FE_OFN484_n4675));
   AO22XLTS U2077 (.Y(n6236), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[29] ), 
	.B0(FE_OFN470_n4676), 
	.A1(FE_OFN1641_acc_fir_data_in_29_), 
	.A0(FE_OFN477_n4675));
   AO22XLTS U2105 (.Y(n6264), 
	.B1(\fifo_from_fir/fifo_cell15/sr_out[1] ), 
	.B0(FE_OFN463_n4676), 
	.A1(FE_OFN1805_acc_fir_data_in_1_), 
	.A0(FE_OFN480_n4675));
   AO22XLTS U1459 (.Y(n5720), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[16] ), 
	.B0(FE_OFN138_n4490), 
	.A1(FE_OFN1533_acc_fft_data_in_16_), 
	.A0(FE_OFN150_n4489));
   AO22XLTS U1475 (.Y(n5736), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[0] ), 
	.B0(FE_OFN132_n4490), 
	.A1(FE_OFN1623_acc_fft_data_in_0_), 
	.A0(FE_OFN144_n4489));
   AO22XLTS U1453 (.Y(n5714), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[22] ), 
	.B0(FE_OFN135_n4490), 
	.A1(FE_OFN1498_acc_fft_data_in_22_), 
	.A0(FE_OFN147_n4489));
   AO22XLTS U1457 (.Y(n5718), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[18] ), 
	.B0(FE_OFN129_n4490), 
	.A1(FE_OFN1525_acc_fft_data_in_18_), 
	.A0(FE_OFN143_n4489));
   AO22XLTS U1473 (.Y(n5734), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[2] ), 
	.B0(FE_OFN133_n4490), 
	.A1(FE_OFN1609_acc_fft_data_in_2_), 
	.A0(FE_OFN141_n4489));
   AO22XLTS U1458 (.Y(n5719), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[17] ), 
	.B0(FE_OFN138_n4490), 
	.A1(FE_OFN1529_acc_fft_data_in_17_), 
	.A0(FE_OFN150_n4489));
   AO22XLTS U1452 (.Y(n5713), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[23] ), 
	.B0(FE_OFN130_n4490), 
	.A1(FE_OFN1496_acc_fft_data_in_23_), 
	.A0(FE_OFN145_n4489));
   AO22XLTS U1474 (.Y(n5735), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[1] ), 
	.B0(FE_OFN133_n4490), 
	.A1(FE_OFN1617_acc_fft_data_in_1_), 
	.A0(FE_OFN141_n4489));
   AO22XLTS U1472 (.Y(n5733), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[3] ), 
	.B0(FE_OFN132_n4490), 
	.A1(FE_OFN1604_acc_fft_data_in_3_), 
	.A0(FE_OFN144_n4489));
   AO22XLTS U1454 (.Y(n5715), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[21] ), 
	.B0(FE_OFN135_n4490), 
	.A1(FE_OFN1509_acc_fft_data_in_21_), 
	.A0(FE_OFN147_n4489));
   AO22XLTS U1456 (.Y(n5717), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[19] ), 
	.B0(FE_OFN129_n4490), 
	.A1(FE_OFN1518_acc_fft_data_in_19_), 
	.A0(FE_OFN143_n4489));
   AO22XLTS U1455 (.Y(n5716), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[20] ), 
	.B0(FE_OFN130_n4490), 
	.A1(FE_OFN1514_acc_fft_data_in_20_), 
	.A0(FE_OFN145_n4489));
   AO22XLTS U1445 (.Y(n5706), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[30] ), 
	.B0(FE_OFN134_n4490), 
	.A1(FE_OFN1460_acc_fft_data_in_30_), 
	.A0(FE_OFN146_n4489));
   AO22XLTS U1448 (.Y(n5709), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[27] ), 
	.B0(FE_OFN131_n4490), 
	.A1(FE_OFN1474_acc_fft_data_in_27_), 
	.A0(FE_OFN141_n4489));
   AO22XLTS U1461 (.Y(n5722), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[14] ), 
	.B0(FE_OFN138_n4490), 
	.A1(FE_OFN1546_acc_fft_data_in_14_), 
	.A0(FE_OFN150_n4489));
   AO22XLTS U1447 (.Y(n5708), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[28] ), 
	.B0(FE_OFN134_n4490), 
	.A1(FE_OFN1472_acc_fft_data_in_28_), 
	.A0(FE_OFN146_n4489));
   AO22XLTS U1466 (.Y(n5727), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[9] ), 
	.B0(FE_OFN136_n4490), 
	.A1(FE_OFN1571_acc_fft_data_in_9_), 
	.A0(FE_OFN148_n4489));
   AO22XLTS U1446 (.Y(n5707), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[29] ), 
	.B0(FE_OFN134_n4490), 
	.A1(FE_OFN1464_acc_fft_data_in_29_), 
	.A0(FE_OFN146_n4489));
   AO22XLTS U1450 (.Y(n5711), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[25] ), 
	.B0(FE_OFN133_n4490), 
	.A1(FE_OFN1484_acc_fft_data_in_25_), 
	.A0(FE_OFN140_n4489));
   AO22XLTS U1462 (.Y(n5723), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[13] ), 
	.B0(FE_OFN137_n4490), 
	.A1(FE_OFN1549_acc_fft_data_in_13_), 
	.A0(FE_OFN149_n4489));
   AO22XLTS U1465 (.Y(n5726), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[10] ), 
	.B0(FE_OFN136_n4490), 
	.A1(FE_OFN1565_acc_fft_data_in_10_), 
	.A0(FE_OFN148_n4489));
   AO22XLTS U1467 (.Y(n5728), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[8] ), 
	.B0(FE_OFN136_n4490), 
	.A1(FE_OFN1579_acc_fft_data_in_8_), 
	.A0(FE_OFN148_n4489));
   AO22XLTS U1451 (.Y(n5712), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[24] ), 
	.B0(FE_OFN133_n4490), 
	.A1(FE_OFN1490_acc_fft_data_in_24_), 
	.A0(FE_OFN140_n4489));
   AO22XLTS U1444 (.Y(n5705), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[31] ), 
	.B0(FE_OFN135_n4490), 
	.A1(FE_OFN1453_acc_fft_data_in_31_), 
	.A0(FE_OFN147_n4489));
   AO22XLTS U1460 (.Y(n5721), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[15] ), 
	.B0(FE_OFN137_n4490), 
	.A1(FE_OFN1542_acc_fft_data_in_15_), 
	.A0(FE_OFN149_n4489));
   AO22XLTS U1464 (.Y(n5725), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[11] ), 
	.B0(FE_OFN137_n4490), 
	.A1(FE_OFN1559_acc_fft_data_in_11_), 
	.A0(FE_OFN149_n4489));
   AO22XLTS U1463 (.Y(n5724), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[12] ), 
	.B0(FE_OFN138_n4490), 
	.A1(FE_OFN1554_acc_fft_data_in_12_), 
	.A0(FE_OFN150_n4489));
   AO22XLTS U1449 (.Y(n5710), 
	.B1(\fifo_from_fft/fifo_cell15/sr_out[26] ), 
	.B0(FE_OFN132_n4490), 
	.A1(FE_OFN1479_acc_fft_data_in_26_), 
	.A0(FE_OFN144_n4489));
   AO22XLTS U749 (.Y(n5429), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[22] ), 
	.B0(FE_OFN70_n3797), 
	.A1(FE_OFN1501_acc_fft_data_in_22_), 
	.A0(FE_OFN80_n3796));
   AO22XLTS U705 (.Y(n5396), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[20] ), 
	.B0(FE_OFN401_n3777), 
	.A1(FE_OFN1692_acc_fir_data_in_20_), 
	.A0(FE_OFN419_n3776));
   AO22XLTS U741 (.Y(n5421), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[30] ), 
	.B0(FE_OFN68_n3797), 
	.A1(FE_OFN1461_acc_fft_data_in_30_), 
	.A0(FE_OFN78_n3796));
   AO22XLTS U754 (.Y(n5434), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[17] ), 
	.B0(FE_OFN71_n3797), 
	.A1(FE_OFN1530_acc_fft_data_in_17_), 
	.A0(FE_OFN83_n3796));
   AO22XLTS U702 (.Y(n5393), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[23] ), 
	.B0(FE_OFN406_n3777), 
	.A1(FE_OFN1671_acc_fir_data_in_23_), 
	.A0(FE_OFN418_n3776));
   AO22XLTS U753 (.Y(n5433), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[18] ), 
	.B0(FE_OFN67_n3797), 
	.A1(FE_OFN1524_acc_fft_data_in_18_), 
	.A0(FE_OFN79_n3796));
   AO22XLTS U755 (.Y(n5435), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[16] ), 
	.B0(FE_OFN71_n3797), 
	.A1(FE_OFN1535_acc_fft_data_in_16_), 
	.A0(FE_OFN83_n3796));
   AO22XLTS U742 (.Y(n5422), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[29] ), 
	.B0(FE_OFN68_n3797), 
	.A1(FE_OFN1466_acc_fft_data_in_29_), 
	.A0(FE_OFN78_n3796));
   AO22XLTS U740 (.Y(n5420), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[31] ), 
	.B0(FE_OFN70_n3797), 
	.A1(FE_OFN1453_acc_fft_data_in_31_), 
	.A0(FE_OFN80_n3796));
   AO22XLTS U748 (.Y(n5428), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[23] ), 
	.B0(FE_OFN65_n3797), 
	.A1(FE_OFN1497_acc_fft_data_in_23_), 
	.A0(FE_OFN77_n3796));
   AO22XLTS U752 (.Y(n5432), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[19] ), 
	.B0(FE_OFN67_n3797), 
	.A1(FE_OFN1516_acc_fft_data_in_19_), 
	.A0(FE_OFN79_n3796));
   AO22XLTS U704 (.Y(n5395), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[21] ), 
	.B0(FE_OFN401_n3777), 
	.A1(FE_OFN1689_acc_fir_data_in_21_), 
	.A0(FE_OFN419_n3776));
   AO22XLTS U703 (.Y(n5394), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[22] ), 
	.B0(FE_OFN401_n3777), 
	.A1(FE_OFN1680_acc_fir_data_in_22_), 
	.A0(FE_OFN422_n3776));
   AO22XLTS U751 (.Y(n5431), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[20] ), 
	.B0(FE_OFN69_n3797), 
	.A1(FE_OFN1510_acc_fft_data_in_20_), 
	.A0(FE_OFN81_n3796));
   AO22XLTS U750 (.Y(n5430), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[21] ), 
	.B0(FE_OFN70_n3797), 
	.A1(FE_OFN1509_acc_fft_data_in_21_), 
	.A0(FE_OFN80_n3796));
   AO22XLTS U706 (.Y(n5397), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[19] ), 
	.B0(FE_OFN406_n3777), 
	.A1(FE_OFN1695_acc_fir_data_in_19_), 
	.A0(FE_OFN416_n3776));
   AO22XLTS U708 (.Y(n5399), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[17] ), 
	.B0(FE_OFN409_n3777), 
	.A1(FE_OFN1709_acc_fir_data_in_17_), 
	.A0(FE_OFN418_n3776));
   AO22XLTS U701 (.Y(n5392), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[24] ), 
	.B0(FE_OFN408_n3777), 
	.A1(FE_OFN1669_acc_fir_data_in_24_), 
	.A0(FE_OFN412_n3776));
   AO22XLTS U719 (.Y(n5410), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[6] ), 
	.B0(FE_OFN404_n3777), 
	.A1(FE_OFN1774_acc_fir_data_in_6_), 
	.A0(FE_OFN415_n3776));
   AO22XLTS U707 (.Y(n5398), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[18] ), 
	.B0(FE_OFN409_n3777), 
	.A1(FE_OFN1704_acc_fir_data_in_18_), 
	.A0(FE_OFN420_n3776));
   AO22XLTS U723 (.Y(n5414), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[2] ), 
	.B0(FE_OFN406_n3777), 
	.A1(FE_OFN1797_acc_fir_data_in_2_), 
	.A0(FE_OFN416_n3776));
   AO22XLTS U721 (.Y(n5412), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[4] ), 
	.B0(FE_OFN402_n3777), 
	.A1(FE_OFN1786_acc_fir_data_in_4_), 
	.A0(FE_OFN415_n3776));
   AO22XLTS U743 (.Y(n5423), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[28] ), 
	.B0(FE_OFN68_n3797), 
	.A1(FE_OFN1472_acc_fft_data_in_28_), 
	.A0(FE_OFN78_n3796));
   AO22XLTS U695 (.Y(n5386), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[30] ), 
	.B0(FE_OFN410_n3777), 
	.A1(FE_OFN1637_acc_fir_data_in_30_), 
	.A0(FE_OFN414_n3776));
   AO22XLTS U697 (.Y(n5388), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[28] ), 
	.B0(FE_OFN410_n3777), 
	.A1(FE_OFN1646_acc_fir_data_in_28_), 
	.A0(FE_OFN414_n3776));
   AO22XLTS U694 (.Y(n5385), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[31] ), 
	.B0(FE_OFN410_n3777), 
	.A1(FE_OFN1632_acc_fir_data_in_31_), 
	.A0(FE_OFN414_n3776));
   AO22XLTS U710 (.Y(n5401), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[15] ), 
	.B0(FE_OFN405_n3777), 
	.A1(FE_OFN1722_acc_fir_data_in_15_), 
	.A0(FE_OFN420_n3776));
   AO22XLTS U717 (.Y(n5408), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[8] ), 
	.B0(FE_OFN411_n3777), 
	.A1(FE_OFN1758_acc_fir_data_in_8_), 
	.A0(FE_OFN421_n3776));
   AO22XLTS U714 (.Y(n5405), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[11] ), 
	.B0(FE_OFN411_n3777), 
	.A1(FE_OFN1741_acc_fir_data_in_11_), 
	.A0(FE_OFN421_n3776));
   AO22XLTS U700 (.Y(n5391), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[25] ), 
	.B0(FE_OFN408_n3777), 
	.A1(FE_OFN1664_acc_fir_data_in_25_), 
	.A0(FE_OFN412_n3776));
   AO22XLTS U712 (.Y(n5403), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[13] ), 
	.B0(FE_OFN411_n3777), 
	.A1(FE_OFN1732_acc_fir_data_in_13_), 
	.A0(FE_OFN421_n3776));
   AO22XLTS U722 (.Y(n5413), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[3] ), 
	.B0(FE_OFN403_n3777), 
	.A1(FE_OFN1793_acc_fir_data_in_3_), 
	.A0(FE_OFN417_n3776));
   AO22XLTS U696 (.Y(n5387), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[29] ), 
	.B0(FE_OFN410_n3777), 
	.A1(FE_OFN1645_acc_fir_data_in_29_), 
	.A0(FE_OFN414_n3776));
   AO22XLTS U709 (.Y(n5400), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[16] ), 
	.B0(FE_OFN409_n3777), 
	.A1(FE_OFN1713_acc_fir_data_in_16_), 
	.A0(FE_OFN418_n3776));
   AO22XLTS U698 (.Y(n5389), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[27] ), 
	.B0(FE_OFN407_n3777), 
	.A1(FE_OFN1655_acc_fir_data_in_27_), 
	.A0(FE_OFN413_n3776));
   AO22XLTS U724 (.Y(n5415), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[1] ), 
	.B0(n3777), 
	.A1(FE_OFN1806_acc_fir_data_in_1_), 
	.A0(FE_OFN419_n3776));
   AO22XLTS U718 (.Y(n5409), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[7] ), 
	.B0(FE_OFN404_n3777), 
	.A1(FE_OFN1767_acc_fir_data_in_7_), 
	.A0(FE_OFN415_n3776));
   AO22XLTS U725 (.Y(n5416), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[0] ), 
	.B0(FE_OFN403_n3777), 
	.A1(FE_OFN1817_acc_fir_data_in_0_), 
	.A0(FE_OFN417_n3776));
   AO22XLTS U716 (.Y(n5407), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[9] ), 
	.B0(FE_OFN411_n3777), 
	.A1(FE_OFN1753_acc_fir_data_in_9_), 
	.A0(FE_OFN421_n3776));
   AO22XLTS U720 (.Y(n5411), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[5] ), 
	.B0(FE_OFN404_n3777), 
	.A1(FE_OFN1781_acc_fir_data_in_5_), 
	.A0(FE_OFN412_n3776));
   AO22XLTS U699 (.Y(n5390), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[26] ), 
	.B0(FE_OFN407_n3777), 
	.A1(FE_OFN1657_acc_fir_data_in_26_), 
	.A0(FE_OFN413_n3776));
   AO22XLTS U715 (.Y(n5406), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[10] ), 
	.B0(FE_OFN405_n3777), 
	.A1(FE_OFN1750_acc_fir_data_in_10_), 
	.A0(FE_OFN422_n3776));
   AO22XLTS U711 (.Y(n5402), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[14] ), 
	.B0(FE_OFN405_n3777), 
	.A1(FE_OFN1729_acc_fir_data_in_14_), 
	.A0(FE_OFN422_n3776));
   AO22XLTS U713 (.Y(n5404), 
	.B1(\fifo_from_fir/fifo_cell0/sr_out[12] ), 
	.B0(FE_OFN405_n3777), 
	.A1(FE_OFN1740_acc_fir_data_in_12_), 
	.A0(FE_OFN422_n3776));
   AO22XLTS U761 (.Y(n5441), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[10] ), 
	.B0(FE_OFN72_n3797), 
	.A1(FE_OFN1568_acc_fft_data_in_10_), 
	.A0(FE_OFN82_n3796));
   AO22XLTS U760 (.Y(n5440), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[11] ), 
	.B0(FE_OFN72_n3797), 
	.A1(FE_OFN1561_acc_fft_data_in_11_), 
	.A0(FE_OFN82_n3796));
   OAI21XLTS U733 (.Y(n3791), 
	.B0(n9489), 
	.A1(n3784), 
	.A0(n3783));
   AO22XLTS U764 (.Y(n5444), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[7] ), 
	.B0(n3797), 
	.A1(FE_OFN1581_acc_fft_data_in_7_), 
	.A0(FE_OFN73_n3796));
   AO22XLTS U769 (.Y(n5449), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[2] ), 
	.B0(FE_OFN63_n3797), 
	.A1(FE_OFN1608_acc_fft_data_in_2_), 
	.A0(FE_OFN74_n3796));
   AO22XLTS U745 (.Y(n5425), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[26] ), 
	.B0(FE_OFN64_n3797), 
	.A1(FE_OFN1478_acc_fft_data_in_26_), 
	.A0(FE_OFN77_n3796));
   AO22XLTS U762 (.Y(n5442), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[9] ), 
	.B0(FE_OFN72_n3797), 
	.A1(FE_OFN1571_acc_fft_data_in_9_), 
	.A0(FE_OFN82_n3796));
   AO22XLTS U763 (.Y(n5443), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[8] ), 
	.B0(FE_OFN72_n3797), 
	.A1(FE_OFN1579_acc_fft_data_in_8_), 
	.A0(FE_OFN82_n3796));
   AO22XLTS U771 (.Y(n5451), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[0] ), 
	.B0(FE_OFN66_n3797), 
	.A1(FE_OFN1623_acc_fft_data_in_0_), 
	.A0(FE_OFN76_n3796));
   AO22XLTS U746 (.Y(n5426), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[25] ), 
	.B0(FE_OFN63_n3797), 
	.A1(FE_OFN1483_acc_fft_data_in_25_), 
	.A0(FE_OFN74_n3796));
   AO22XLTS U757 (.Y(n5437), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[14] ), 
	.B0(FE_OFN71_n3797), 
	.A1(FE_OFN1546_acc_fft_data_in_14_), 
	.A0(FE_OFN83_n3796));
   AO22XLTS U758 (.Y(n5438), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[13] ), 
	.B0(FE_OFN69_n3797), 
	.A1(FE_OFN1550_acc_fft_data_in_13_), 
	.A0(FE_OFN81_n3796));
   AO22XLTS U744 (.Y(n5424), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[27] ), 
	.B0(FE_OFN66_n3797), 
	.A1(FE_OFN1473_acc_fft_data_in_27_), 
	.A0(FE_OFN75_n3796));
   AO22XLTS U765 (.Y(n5445), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[6] ), 
	.B0(FE_OFN67_n3797), 
	.A1(FE_OFN1586_acc_fft_data_in_6_), 
	.A0(FE_OFN79_n3796));
   AO22XLTS U770 (.Y(n5450), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[1] ), 
	.B0(FE_OFN64_n3797), 
	.A1(FE_OFN1615_acc_fft_data_in_1_), 
	.A0(FE_OFN75_n3796));
   AO22XLTS U747 (.Y(n5427), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[24] ), 
	.B0(FE_OFN63_n3797), 
	.A1(FE_OFN1490_acc_fft_data_in_24_), 
	.A0(FE_OFN74_n3796));
   AO22XLTS U768 (.Y(n5448), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[3] ), 
	.B0(FE_OFN66_n3797), 
	.A1(FE_OFN1604_acc_fft_data_in_3_), 
	.A0(FE_OFN76_n3796));
   AO22XLTS U756 (.Y(n5436), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[15] ), 
	.B0(FE_OFN69_n3797), 
	.A1(FE_OFN1542_acc_fft_data_in_15_), 
	.A0(FE_OFN81_n3796));
   AO22XLTS U766 (.Y(n5446), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[5] ), 
	.B0(FE_OFN65_n3797), 
	.A1(FE_OFN1594_acc_fft_data_in_5_), 
	.A0(FE_OFN77_n3796));
   AO22XLTS U759 (.Y(n5439), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[12] ), 
	.B0(FE_OFN71_n3797), 
	.A1(FE_OFN1556_acc_fft_data_in_12_), 
	.A0(FE_OFN83_n3796));
   AO22XLTS U767 (.Y(n5447), 
	.B1(\fifo_from_fft/fifo_cell0/sr_out[4] ), 
	.B0(n3797), 
	.A1(FE_OFN1598_acc_fft_data_in_4_), 
	.A0(FE_OFN73_n3796));
   OAI21XLTS U687 (.Y(n3771), 
	.B0(n9488), 
	.A1(n3764), 
	.A0(n3763));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[25]  (.QN(\router/addr_calc/iir_read_calc/count[25] ), 
	.Q(n8020), 
	.D(n7087), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[24]  (.QN(\router/addr_calc/iir_read_calc/count[24] ), 
	.Q(n8031), 
	.D(n7086), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[23]  (.QN(\router/addr_calc/iir_read_calc/count[23] ), 
	.Q(n8021), 
	.D(n7085), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[22]  (.QN(\router/addr_calc/iir_read_calc/count[22] ), 
	.Q(n8032), 
	.D(n7084), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[29]  (.QN(\router/addr_calc/iir_read_calc/count[29] ), 
	.Q(n8012), 
	.D(n7083), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[28]  (.QN(\router/addr_calc/iir_read_calc/count[28] ), 
	.Q(n8016), 
	.D(n7082), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[27]  (.QN(\router/addr_calc/iir_read_calc/count[27] ), 
	.Q(n8019), 
	.D(n7081), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[26]  (.QN(\router/addr_calc/iir_read_calc/count[26] ), 
	.Q(n8030), 
	.D(n7080), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[21]  (.QN(\router/addr_calc/iir_read_calc/count[21] ), 
	.Q(n8022), 
	.D(n7079), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[20]  (.QN(\router/addr_calc/iir_read_calc/count[20] ), 
	.Q(n8033), 
	.D(n7078), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[19]  (.QN(\router/addr_calc/iir_read_calc/count[19] ), 
	.Q(n8023), 
	.D(n7077), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[18]  (.QN(\router/addr_calc/iir_read_calc/count[18] ), 
	.Q(n8034), 
	.D(n7076), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[31]  (.QN(\router/addr_calc/iir_read_calc/count[31] ), 
	.Q(n8014), 
	.D(n7075), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[10]  (.QN(\router/addr_calc/iir_read_calc/count[10] ), 
	.Q(n8038), 
	.D(n7074), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[9]  (.QN(\router/addr_calc/iir_read_calc/count[9] ), 
	.Q(n8028), 
	.D(n7073), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[8]  (.QN(\router/addr_calc/iir_read_calc/count[8] ), 
	.Q(n8039), 
	.D(n7072), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[7]  (.QN(\router/addr_calc/iir_read_calc/count[7] ), 
	.Q(n8029), 
	.D(n7071), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[6]  (.QN(\router/addr_calc/iir_read_calc/count[6] ), 
	.Q(n8040), 
	.D(n7070), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[5]  (.QN(\router/addr_calc/iir_read_calc/count[5] ), 
	.Q(n8013), 
	.D(n7069), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[4]  (.QN(\router/addr_calc/iir_read_calc/count[4] ), 
	.Q(n8017), 
	.D(n7068), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[3]  (.QN(\router/addr_calc/iir_read_calc/count[3] ), 
	.Q(n8041), 
	.D(n7067), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[2]  (.QN(\router/addr_calc/iir_read_calc/count[2] ), 
	.Q(n8042), 
	.D(n7066), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[1]  (.QN(\router/addr_calc/iir_read_calc/count[1] ), 
	.Q(n8015), 
	.D(n7065), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[0]  (.QN(\router/addr_calc/iir_read_calc/count[0] ), 
	.Q(n8018), 
	.D(n7064), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[30]  (.QN(\router/addr_calc/iir_read_calc/count[30] ), 
	.Q(n8011), 
	.D(n7063), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[17]  (.QN(\router/addr_calc/iir_read_calc/count[17] ), 
	.Q(n8024), 
	.D(n7062), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[16]  (.QN(\router/addr_calc/iir_read_calc/count[16] ), 
	.Q(n8035), 
	.D(n7061), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[15]  (.QN(\router/addr_calc/iir_read_calc/count[15] ), 
	.Q(n8025), 
	.D(n7060), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[14]  (.QN(\router/addr_calc/iir_read_calc/count[14] ), 
	.Q(n8036), 
	.D(n7059), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[13]  (.QN(\router/addr_calc/iir_read_calc/count[13] ), 
	.Q(n8026), 
	.D(n7058), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[12]  (.QN(\router/addr_calc/iir_read_calc/count[12] ), 
	.Q(n8037), 
	.D(n7057), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/iir_read_calc/counter/count_reg[11]  (.QN(\router/addr_calc/iir_read_calc/count[11] ), 
	.Q(n8027), 
	.D(n7056), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[2]  (.QN(n7106), 
	.Q(n7107), 
	.E(FE_OFN1199_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N180 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[1]  (.QN(n7111), 
	.Q(n7112), 
	.E(n7014), 
	.D(\router/addr_calc/iir_write_calc/counter/N179 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[7]  (.QN(n7091), 
	.Q(n7093), 
	.E(FE_OFN1207_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N185 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[6]  (.QN(n7088), 
	.Q(n7090), 
	.E(FE_OFN1207_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N184 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[5]  (.Q(\router/addr_calc/iir_write_calc/count[5] ), 
	.E(n7014), 
	.D(\router/addr_calc/iir_write_calc/counter/N183 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[4]  (.QN(n7094), 
	.Q(n7095), 
	.E(FE_OFN1199_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N182 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[8]  (.QN(n7097), 
	.Q(n7099), 
	.E(FE_OFN1204_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N186 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[3]  (.QN(n7100), 
	.Q(n7102), 
	.E(FE_OFN1207_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N181 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[9]  (.Q(\router/addr_calc/iir_write_calc/count[9] ), 
	.E(FE_OFN1206_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N187 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[10]  (.QN(n7103), 
	.Q(n7105), 
	.E(FE_OFN1206_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N188 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[11]  (.QN(n7108), 
	.Q(n7110), 
	.E(FE_OFN1204_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N189 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[12]  (.QN(n7114), 
	.Q(n7116), 
	.E(FE_OFN1203_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N190 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[13]  (.QN(n7120), 
	.Q(n7122), 
	.E(FE_OFN1205_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N191 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[14]  (.QN(n7125), 
	.Q(n7127), 
	.E(FE_OFN1205_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N192 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[10]  (.QN(n7327), 
	.Q(n7328), 
	.E(FE_OFN1193_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N188 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[8]  (.QN(n7332), 
	.Q(n7333), 
	.E(FE_OFN1192_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N186 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[10]  (.QN(n7441), 
	.Q(n7443), 
	.E(FE_OFN1162_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N188 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[8]  (.QN(n7446), 
	.Q(n7448), 
	.E(FE_OFN1161_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N186 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[1]  (.QN(n7362), 
	.Q(n7363), 
	.E(FE_OFN1191_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N179 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[10]  (.QN(n7565), 
	.Q(n7567), 
	.E(FE_OFN1175_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N188 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[8]  (.QN(n7570), 
	.Q(n7572), 
	.E(FE_OFN1175_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N186 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[14]  (.QN(n7307), 
	.Q(n7308), 
	.E(FE_OFN1194_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N192 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[13]  (.QN(n7312), 
	.Q(n7314), 
	.E(FE_OFN1193_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N191 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[12]  (.QN(n7317), 
	.Q(n7319), 
	.E(FE_OFN1194_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N190 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[7]  (.QN(n7337), 
	.Q(n7339), 
	.E(FE_OFN1192_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N185 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[6]  (.QN(n7342), 
	.Q(n7344), 
	.E(FE_OFN1192_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N184 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[5]  (.Q(\router/addr_calc/fir_read_calc/count[5] ), 
	.E(n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N183 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[4]  (.QN(n7347), 
	.Q(n7348), 
	.E(FE_OFN1191_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N182 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[3]  (.QN(n7352), 
	.Q(n7353), 
	.E(FE_OFN1190_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N181 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[2]  (.QN(n7357), 
	.Q(n7358), 
	.E(n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N180 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[14]  (.QN(n7421), 
	.Q(n7423), 
	.E(FE_OFN1167_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N192 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[13]  (.QN(n7426), 
	.Q(n7428), 
	.E(FE_OFN1164_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N191 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[12]  (.QN(n7431), 
	.Q(n7433), 
	.E(FE_OFN1164_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N190 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[7]  (.QN(n7451), 
	.Q(n7453), 
	.E(FE_OFN1161_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N185 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[1]  (.QN(n7481), 
	.Q(n7482), 
	.E(FE_OFN1159_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N179 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[5]  (.QN(n7461), 
	.Q(n7462), 
	.E(n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N183 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[4]  (.QN(n7466), 
	.Q(n7467), 
	.E(FE_OFN1158_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N182 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[6]  (.QN(n7456), 
	.Q(n7458), 
	.E(FE_OFN1158_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N184 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[3]  (.QN(n7471), 
	.Q(n7473), 
	.E(n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N181 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[2]  (.QN(n7476), 
	.Q(n7478), 
	.E(FE_OFN1158_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N180 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[1]  (.QN(n7600), 
	.Q(n7601), 
	.E(FE_OFN1170_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N179 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[5]  (.Q(\router/addr_calc/fft_read_calc/count[5] ), 
	.E(FE_OFN1174_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N183 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[4]  (.QN(n7585), 
	.Q(n7586), 
	.E(FE_OFN1176_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N182 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[14]  (.QN(n7545), 
	.Q(n7547), 
	.E(FE_OFN1178_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N192 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[13]  (.QN(n7550), 
	.Q(n7552), 
	.E(FE_OFN1177_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N191 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[12]  (.QN(n7555), 
	.Q(n7557), 
	.E(FE_OFN1178_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N190 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[7]  (.QN(n7575), 
	.Q(n7577), 
	.E(FE_OFN1178_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N185 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[6]  (.QN(n7580), 
	.Q(n7582), 
	.E(FE_OFN1176_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N184 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[3]  (.QN(n7590), 
	.Q(n7592), 
	.E(FE_OFN1169_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N181 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[2]  (.QN(n7595), 
	.Q(n7597), 
	.E(FE_OFN1169_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N180 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[10]  (.QN(n7208), 
	.Q(n7210), 
	.E(FE_OFN1185_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N188 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[8]  (.QN(n7213), 
	.Q(n7215), 
	.E(FE_OFN1185_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N186 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[1]  (.QN(n7243), 
	.Q(n7244), 
	.E(FE_OFN1188_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N179 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[14]  (.QN(n7188), 
	.Q(n7190), 
	.E(FE_OFN1189_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N192 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[13]  (.QN(n7194), 
	.Q(n7196), 
	.E(FE_OFN1186_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N191 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[4]  (.QN(n7228), 
	.Q(n7229), 
	.E(FE_OFN1182_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N182 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[3]  (.QN(n7233), 
	.Q(n7235), 
	.E(FE_OFN1181_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N181 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[2]  (.QN(n7238), 
	.Q(n7240), 
	.E(FE_OFN1187_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N180 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[12]  (.QN(n7200), 
	.Q(n7202), 
	.E(FE_OFN1186_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N190 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[5]  (.Q(\router/addr_calc/fir_write_calc/count[5] ), 
	.E(FE_OFN1180_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N183 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[7]  (.QN(n7218), 
	.Q(n7220), 
	.E(FE_OFN1182_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N185 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[6]  (.QN(n7223), 
	.Q(n7225), 
	.E(FE_OFN1182_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N184 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[15]  (.QN(n7182), 
	.Q(n7184), 
	.E(FE_OFN1189_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N193 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[15]  (.Q(\router/addr_calc/fir_read_calc/count[15] ), 
	.E(FE_OFN1193_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N193 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[15]  (.Q(\router/addr_calc/fft_write_calc/count[15] ), 
	.E(FE_OFN1164_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N193 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[15]  (.QN(n7540), 
	.Q(n7542), 
	.E(FE_OFN1177_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N193 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[11]  (.QN(n7322), 
	.Q(n7323), 
	.E(FE_OFN1192_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N189 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[9]  (.Q(\router/addr_calc/fir_read_calc/count[9] ), 
	.E(n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N187 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[11]  (.QN(n7436), 
	.Q(n7438), 
	.E(FE_OFN1162_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N189 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[9]  (.Q(\router/addr_calc/fft_write_calc/count[9] ), 
	.E(FE_OFN1162_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N187 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[11]  (.QN(n7560), 
	.Q(n7562), 
	.E(FE_OFN1175_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N189 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[9]  (.Q(\router/addr_calc/fft_read_calc/count[9] ), 
	.E(FE_OFN1178_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N187 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[15]  (.QN(n7131), 
	.Q(n7133), 
	.E(FE_OFN1203_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N193 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[11]  (.QN(n7204), 
	.Q(n7206), 
	.E(FE_OFN1186_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N189 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[9]  (.Q(\router/addr_calc/fir_write_calc/count[9] ), 
	.E(FE_OFN1185_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N187 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[16]  (.QN(n7302), 
	.Q(n7303), 
	.E(FE_OFN1194_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N194 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[16]  (.Q(\router/addr_calc/fir_write_calc/count[16] ), 
	.E(FE_OFN1189_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N194 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[16]  (.Q(\router/addr_calc/fft_read_calc/count[16] ), 
	.E(FE_OFN1177_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N194 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[16]  (.QN(n7416), 
	.Q(n7418), 
	.E(FE_OFN1167_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N194 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[17]  (.QN(n7176), 
	.Q(n7178), 
	.E(FE_OFN1188_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N195 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[17]  (.QN(n7297), 
	.Q(n7298), 
	.E(FE_OFN1195_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N195 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[17]  (.QN(n7411), 
	.Q(n7413), 
	.E(FE_OFN1167_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N195 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[17]  (.QN(n7535), 
	.Q(n7537), 
	.E(FE_OFN1177_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N195 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[17]  (.QN(n7137), 
	.Q(n7139), 
	.E(FE_OFN1205_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N195 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[18]  (.QN(n7170), 
	.Q(n7171), 
	.E(FE_OFN1188_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N196 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[18]  (.QN(n7292), 
	.Q(n7293), 
	.E(FE_OFN1195_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N196 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[18]  (.QN(n7406), 
	.Q(n7407), 
	.E(FE_OFN1165_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N196 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[18]  (.QN(n7530), 
	.Q(n7531), 
	.E(FE_OFN1173_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N196 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[18]  (.QN(n7143), 
	.Q(n7144), 
	.E(FE_OFN1202_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N196 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[19]  (.Q(\router/addr_calc/fir_write_calc/count[19] ), 
	.E(FE_OFN1189_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N197 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[19]  (.Q(\router/addr_calc/fir_read_calc/count[19] ), 
	.E(FE_OFN1198_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N197 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[19]  (.Q(\router/addr_calc/fft_write_calc/count[19] ), 
	.E(FE_OFN1165_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N197 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[19]  (.Q(\router/addr_calc/fft_read_calc/count[19] ), 
	.E(FE_OFN1173_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N197 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[20]  (.QN(n7149), 
	.Q(n7150), 
	.E(FE_OFN1202_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N198 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[20]  (.QN(n7525), 
	.Q(n7526), 
	.E(FE_OFN1173_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N198 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[20]  (.QN(n7164), 
	.Q(n7165), 
	.E(FE_OFN1188_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N198 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[20]  (.QN(n7287), 
	.Q(n7288), 
	.E(FE_OFN1196_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N198 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[20]  (.QN(n7401), 
	.Q(n7402), 
	.E(FE_OFN1165_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N198 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[21]  (.QN(n7158), 
	.Q(n7159), 
	.E(FE_OFN1184_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N199 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[21]  (.QN(n7282), 
	.Q(n7283), 
	.E(FE_OFN1198_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N199 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[21]  (.QN(n7396), 
	.Q(n7397), 
	.E(FE_OFN1165_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N199 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[21]  (.QN(n7520), 
	.Q(n7521), 
	.E(FE_OFN1173_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N199 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[21]  (.QN(n7155), 
	.Q(n7156), 
	.E(FE_OFN1200_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N199 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[22]  (.QN(n7161), 
	.Q(n7163), 
	.E(FE_OFN1200_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N200 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[22]  (.QN(n7515), 
	.Q(n7516), 
	.E(FE_OFN1172_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N200 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[22]  (.QN(n7152), 
	.Q(n7153), 
	.E(FE_OFN1187_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N200 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[22]  (.QN(n7277), 
	.Q(n7278), 
	.E(FE_OFN1196_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N200 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[22]  (.QN(n7391), 
	.Q(n7392), 
	.E(FE_OFN1160_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N200 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[23]  (.Q(\router/addr_calc/fir_write_calc/count[23] ), 
	.E(FE_OFN1184_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N201 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[23]  (.Q(\router/addr_calc/fir_read_calc/count[23] ), 
	.E(FE_OFN1198_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N201 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[23]  (.Q(\router/addr_calc/fft_write_calc/count[23] ), 
	.E(FE_OFN1163_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N201 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[23]  (.Q(\router/addr_calc/fft_read_calc/count[23] ), 
	.E(FE_OFN1171_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N201 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[23]  (.Q(\router/addr_calc/iir_write_calc/count[23] ), 
	.E(FE_OFN1201_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N201 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[24]  (.QN(n7146), 
	.Q(n7148), 
	.E(FE_OFN1184_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N202 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[24]  (.QN(n7272), 
	.Q(n7273), 
	.E(FE_OFN1198_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N202 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[24]  (.QN(n7386), 
	.Q(n7388), 
	.E(FE_OFN1160_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N202 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[24]  (.QN(n7510), 
	.Q(n7512), 
	.E(FE_OFN1171_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N202 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[24]  (.QN(n7167), 
	.Q(n7169), 
	.E(FE_OFN1201_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N202 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[25]  (.QN(n7140), 
	.Q(n7142), 
	.E(FE_OFN1183_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N203 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[25]  (.QN(n7267), 
	.Q(n7268), 
	.E(FE_OFN1196_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N203 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[25]  (.QN(n7381), 
	.Q(n7383), 
	.E(FE_OFN1163_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N203 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[25]  (.QN(n7505), 
	.Q(n7507), 
	.E(FE_OFN1172_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N203 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[25]  (.QN(n7173), 
	.Q(n7175), 
	.E(FE_OFN1204_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N203 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[26]  (.QN(n7134), 
	.Q(n7135), 
	.E(FE_OFN1183_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N204 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[26]  (.QN(n7262), 
	.Q(n7264), 
	.E(FE_OFN1197_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N204 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[26]  (.QN(n7376), 
	.Q(n7377), 
	.E(FE_OFN1166_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N204 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[26]  (.QN(n7500), 
	.Q(n7501), 
	.E(FE_OFN1174_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N204 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[26]  (.QN(n7179), 
	.Q(n7181), 
	.E(FE_OFN1200_router_addr_calc_iir_write_calc_counter_N212), 
	.D(\router/addr_calc/iir_write_calc/counter/N204 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[27]  (.Q(\router/addr_calc/fir_write_calc/count[27] ), 
	.E(FE_OFN1181_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N205 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[27]  (.Q(\router/addr_calc/fir_read_calc/count[27] ), 
	.E(FE_OFN1191_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N205 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[27]  (.Q(\router/addr_calc/fft_write_calc/count[27] ), 
	.E(FE_OFN1166_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N205 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[27]  (.Q(\router/addr_calc/fft_read_calc/count[27] ), 
	.E(FE_OFN1171_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N205 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[28]  (.QN(n7128), 
	.Q(n7129), 
	.E(FE_OFN1181_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N206 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[28]  (.QN(n7257), 
	.Q(n7259), 
	.E(FE_OFN1197_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N206 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[28]  (.QN(n7371), 
	.Q(n7372), 
	.E(FE_OFN1160_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N206 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[28]  (.QN(n7495), 
	.Q(n7496), 
	.E(FE_OFN1170_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N206 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[28]  (.QN(n7185), 
	.Q(n7187), 
	.E(\router/addr_calc/iir_write_calc/counter/N212 ), 
	.D(\router/addr_calc/iir_write_calc/counter/N206 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[29]  (.QN(n7123), 
	.Q(n7124), 
	.E(FE_OFN1179_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N207 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[29]  (.QN(n7253), 
	.Q(n7254), 
	.E(FE_OFN1197_n7023), 
	.D(\router/addr_calc/fir_read_calc/counter/N207 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[29]  (.QN(n7491), 
	.Q(n7492), 
	.E(FE_OFN1168_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N207 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[29]  (.QN(n7191), 
	.Q(n7193), 
	.E(\router/addr_calc/iir_write_calc/counter/N212 ), 
	.D(\router/addr_calc/iir_write_calc/counter/N207 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[29]  (.Q(\router/addr_calc/fft_write_calc/count[29] ), 
	.E(FE_OFN1166_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N207 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[30]  (.QN(n7367), 
	.Q(n7368), 
	.E(FE_OFN1159_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N208 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[30]  (.Q(\router/addr_calc/fir_write_calc/count[30] ), 
	.E(FE_OFN1179_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N208 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[30]  (.Q(\router/addr_calc/fir_read_calc/count[30] ), 
	.E(n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N208 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[30]  (.Q(\router/addr_calc/fft_read_calc/count[30] ), 
	.E(FE_OFN1168_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N208 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_write_calc/counter/count_reg[31]  (.Q(\router/addr_calc/fft_write_calc/count[31] ), 
	.E(FE_OFN1166_n7019), 
	.D(\router/addr_calc/fft_write_calc/counter/N209 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/iir_write_calc/counter/count_reg[31]  (.QN(n7197), 
	.Q(n7198), 
	.E(n7014), 
	.D(\router/addr_calc/iir_write_calc/counter/N209 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_read_calc/counter/count_reg[31]  (.QN(n7248), 
	.Q(n7249), 
	.E(FE_OFN1191_n7022), 
	.D(\router/addr_calc/fir_read_calc/counter/N209 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fir_write_calc/counter/count_reg[31]  (.QN(n7117), 
	.Q(n7118), 
	.E(FE_OFN1180_n7020), 
	.D(\router/addr_calc/fir_write_calc/counter/N209 ), 
	.CK(clk__L1_N0));
   EDFFXLTS \router/addr_calc/fft_read_calc/counter/count_reg[31]  (.QN(n7486), 
	.Q(n7487), 
	.E(FE_OFN1176_n7021), 
	.D(\router/addr_calc/fft_read_calc/counter/N209 ), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/from_fft_go_reg  (.QN(\router/addr_calc/N63 ), 
	.Q(n8063), 
	.D(n5462), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/to_fft_go_reg  (.QN(\router/addr_calc/N9 ), 
	.Q(n8064), 
	.D(n5463), 
	.CK(clk__L1_N0));
   DFFXLTS \fifo_from_fir/empty_det/result_reg  (.QN(n3467), 
	.Q(from_fir_empty), 
	.D(\fifo_from_fir/empty_det/N4 ), 
	.CK(clk__L1_N0));
   DFFXLTS \fifo_from_fft/empty_det/result_reg  (.QN(n3478), 
	.Q(from_fft_empty), 
	.D(\fifo_from_fft/empty_det/N4 ), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/from_fir_go_reg  (.QN(\router/addr_calc/N99 ), 
	.Q(n8061), 
	.D(n5465), 
	.CK(clk__L1_N0));
   DFFXLTS \router/addr_calc/to_fir_go_reg  (.QN(\router/addr_calc/N95 ), 
	.Q(n8062), 
	.D(n5464), 
	.CK(clk__L1_N0));
   DFFXLTS \fifo_to_fir/fifo_cell0/reg_ptok/out_valid_put_reg  (.QN(n3800), 
	.Q(\fifo_to_fir/fifo_cell0/reg_ptok/out_valid_put ), 
	.D(n5453), 
	.CK(clk__L1_N0));
   DFFXLTS \fifo_to_fft/fifo_cell0/reg_ptok/out_valid_put_reg  (.QN(n3811), 
	.Q(\fifo_to_fft/fifo_cell0/reg_ptok/out_valid_put ), 
	.D(n5455), 
	.CK(clk__L1_N0));
   DFFXLTS \fifo_from_fir/fifo_cell0/reg_ptok/out_valid_put_reg  (.QN(n3760), 
	.Q(\fifo_from_fir/fifo_cell0/reg_ptok/out_valid_put ), 
	.D(n5383), 
	.CK(clk__L1_N0));
   DFFXLTS \fifo_from_fft/fifo_cell0/reg_ptok/out_valid_put_reg  (.QN(n3780), 
	.Q(\fifo_from_fft/fifo_cell0/reg_ptok/out_valid_put ), 
	.D(n5418), 
	.CK(clk__L1_N0));
   SDFFQXLTS \router/addr_calc/iir_read_calc/counter/done_reg  (.SI(1'b1), 
	.SE(n9390), 
	.Q(n3710), 
	.D(\router/addr_calc/iir_read_calc/counter/N40 ), 
	.CK(clk__L1_N0));
   OR3X1TS U3895 (.Y(n8055), 
	.C(n4794), 
	.B(n4793), 
	.A(n8872));
   INVX2TS U3898 (.Y(n8784), 
	.A(n8057));
   INVX2TS U3899 (.Y(n8805), 
	.A(FE_OFN730_n8058));
   OR3X1TS U3900 (.Y(n4112), 
	.C(n4170), 
	.B(n4169), 
	.A(n8784));
   OR3X1TS U3901 (.Y(n3937), 
	.C(n3995), 
	.B(n3994), 
	.A(n8805));
   INVX2TS U3902 (.Y(n8785), 
	.A(FE_OFN734_n8057));
   INVX2TS U3903 (.Y(n8806), 
	.A(FE_OFN731_n8058));
   OR3X1TS U3904 (.Y(n4097), 
	.C(n4161), 
	.B(n4160), 
	.A(n8785));
   OR3X1TS U3905 (.Y(n3922), 
	.C(n3986), 
	.B(n3985), 
	.A(n8806));
   INVX2TS U3906 (.Y(n8786), 
	.A(FE_OFN734_n8057));
   OR3X1TS U3907 (.Y(n4092), 
	.C(n4158), 
	.B(n4157), 
	.A(n8785));
   INVX2TS U3908 (.Y(n8807), 
	.A(FE_OFN731_n8058));
   OR3X1TS U3909 (.Y(n3917), 
	.C(n3983), 
	.B(n3982), 
	.A(n8806));
   OR3X1TS U3910 (.Y(n4072), 
	.C(n4146), 
	.B(n4145), 
	.A(n8786));
   OR3X1TS U3911 (.Y(n4077), 
	.C(n4149), 
	.B(n4148), 
	.A(n8786));
   OR3X1TS U3912 (.Y(n3897), 
	.C(n3971), 
	.B(n3970), 
	.A(n8807));
   OR3X1TS U3913 (.Y(n3902), 
	.C(n3974), 
	.B(n3973), 
	.A(n8807));
   NOR3X1TS U3914 (.Y(n3907), 
	.C(n3977), 
	.B(n3976), 
	.A(n8807));
   NOR3X1TS U3915 (.Y(n3932), 
	.C(n3992), 
	.B(n3991), 
	.A(n8806));
   NOR3X1TS U3916 (.Y(n3892), 
	.C(n3968), 
	.B(n3967), 
	.A(n8808));
   NOR3X1TS U3917 (.Y(n4082), 
	.C(n4152), 
	.B(n4151), 
	.A(n8786));
   NOR3X1TS U3918 (.Y(n4107), 
	.C(n4167), 
	.B(n4166), 
	.A(n8785));
   NOR3X1TS U3919 (.Y(n4067), 
	.C(n4143), 
	.B(n4142), 
	.A(n8787));
   NOR3X1TS U3923 (.Y(n4062), 
	.C(n4140), 
	.B(n4139), 
	.A(n8787));
   NOR3X1TS U3924 (.Y(n3887), 
	.C(n3965), 
	.B(n3964), 
	.A(n8808));
   OR2X2TS U3926 (.Y(n7972), 
	.B(FE_OFN700_n3959), 
	.A(FE_OFN797_n7619));
   OR3X1TS U3929 (.Y(n8054), 
	.C(n4608), 
	.B(n4607), 
	.A(n8839));
   OR3X1TS U3944 (.Y(n8053), 
	.C(n4827), 
	.B(n4826), 
	.A(n8870));
   AOI21X1TS U3945 (.Y(n3772), 
	.B0(n3764), 
	.A1(n4674), 
	.A0(\fifo_from_fir/hang[14] ));
   AOI2BB1X1TS U3949 (.Y(n4181), 
	.B0(n3804), 
	.A1N(n4055), 
	.A0N(n4184));
   AOI2BB1X1TS U3951 (.Y(n4006), 
	.B0(n3815), 
	.A1N(n3880), 
	.A0N(n4009));
   ADDHXLTS U3984 (.S(\router/addr_calc/fft_read_calc/counter/N76 ), 
	.CO(\add_x_22_0/carry[31] ), 
	.B(\add_x_22_0/carry[30] ), 
	.A(FE_OFN1229_router_addr_calc_fft_read_calc_count_30_));
   ADDHXLTS U3985 (.S(\router/addr_calc/fir_read_calc/counter/N76 ), 
	.CO(\add_x_22_2/carry[31] ), 
	.B(\add_x_22_2/carry[30] ), 
	.A(FE_OFN1230_router_addr_calc_fir_read_calc_count_30_));
   ADDHXLTS U3986 (.S(\router/addr_calc/fir_write_calc/counter/N76 ), 
	.CO(\add_x_22_3/carry[31] ), 
	.B(\add_x_22_3/carry[30] ), 
	.A(\router/addr_calc/fir_write_calc/count[30] ));
   ADDHXLTS U3987 (.S(\router/addr_calc/iir_write_calc/counter/N75 ), 
	.CO(\add_x_22_5/carry[30] ), 
	.B(\add_x_22_5/carry[29] ), 
	.A(n7193));
   ADDHXLTS U3988 (.S(\router/addr_calc/iir_write_calc/counter/N74 ), 
	.CO(\add_x_22_5/carry[29] ), 
	.B(\add_x_22_5/carry[28] ), 
	.A(n7187));
   ADDHXLTS U3989 (.S(\router/addr_calc/fft_read_calc/counter/N74 ), 
	.CO(\add_x_22_0/carry[29] ), 
	.B(\add_x_22_0/carry[28] ), 
	.A(n7497));
   ADDHXLTS U3992 (.S(\router/addr_calc/fft_write_calc/counter/N74 ), 
	.CO(\add_x_22_1/carry[29] ), 
	.B(\add_x_22_1/carry[28] ), 
	.A(n7373));
   ADDHXLTS U3995 (.S(\router/addr_calc/fir_read_calc/counter/N74 ), 
	.CO(\add_x_22_2/carry[29] ), 
	.B(\add_x_22_2/carry[28] ), 
	.A(FE_OFN1236_n7259));
   ADDHXLTS U3998 (.S(\router/addr_calc/fir_write_calc/counter/N74 ), 
	.CO(\add_x_22_3/carry[29] ), 
	.B(\add_x_22_3/carry[28] ), 
	.A(n7130));
   INVX2TS U4020 (.Y(n9412), 
	.A(FE_OFN989_n9431));
   INVX2TS U4027 (.Y(n9411), 
	.A(FE_OFN989_n9431));
   NAND2X1TS U4032 (.Y(n3530), 
	.B(\router/addr_calc/fir_write_calc/counter/N40 ), 
	.A(\router/data_from_fir ));
   NAND2X1TS U4033 (.Y(n3662), 
	.B(\router/addr_calc/fft_read_calc/counter/N40 ), 
	.A(\router/data_to_fft ));
   NAND2X1TS U4034 (.Y(n3618), 
	.B(\router/addr_calc/fft_write_calc/counter/N40 ), 
	.A(FE_OFN1438_router_data_from_fft));
   NAND2X1TS U4035 (.Y(n3574), 
	.B(\router/addr_calc/fir_read_calc/counter/N40 ), 
	.A(\router/data_to_fir ));
   ADDHXLTS U4044 (.S(\router/addr_calc/fir_write_calc/counter/N47 ), 
	.CO(\add_x_22_3/carry[2] ), 
	.B(FE_OFN1445_router_addr_calc_fir_write_calc_count_0_), 
	.A(n7244));
   ADDHXLTS U4050 (.S(\router/addr_calc/fft_read_calc/counter/N47 ), 
	.CO(\add_x_22_0/carry[2] ), 
	.B(FE_OFN1444_router_addr_calc_fft_read_calc_count_0_), 
	.A(n7601));
   ADDHXLTS U4052 (.S(\router/addr_calc/fft_write_calc/counter/N47 ), 
	.CO(\add_x_22_1/carry[2] ), 
	.B(FE_OFN1443_router_addr_calc_fft_write_calc_count_0_), 
	.A(n7482));
   ADDHXLTS U4061 (.S(\router/addr_calc/fir_read_calc/counter/N47 ), 
	.CO(\add_x_22_2/carry[2] ), 
	.B(\router/addr_calc/fir_read_calc/count[0] ), 
	.A(n7363));
   INVX2TS U4062 (.Y(n9408), 
	.A(FE_OFN985_n9431));
   INVX2TS U4064 (.Y(n9409), 
	.A(FE_OFN989_n9431));
   INVX2TS U4066 (.Y(n9410), 
	.A(FE_OFN987_n9431));
   INVX2TS U4076 (.Y(n9384), 
	.A(FE_OFN1289_iir_enable));
   INVX2TS U4077 (.Y(n9385), 
	.A(FE_OFN1289_iir_enable));
   INVX2TS U4078 (.Y(n9382), 
	.A(FE_OFN1287_iir_enable));
   INVX2TS U4079 (.Y(n9383), 
	.A(FE_OFN1288_iir_enable));
   INVX2TS U4080 (.Y(n9381), 
	.A(FE_OFN1287_iir_enable));
   INVX2TS U4081 (.Y(n9386), 
	.A(FE_OFN1289_iir_enable));
   INVX2TS U4082 (.Y(n9388), 
	.A(FE_OFN1287_iir_enable));
   INVX2TS U4083 (.Y(n9387), 
	.A(FE_OFN1289_iir_enable));
   INVX2TS U4090 (.Y(n4207), 
	.A(n3456));
   INVX2TS U4093 (.Y(n9513), 
	.A(FE_OFN821_n7619));
   NAND2X1TS U4096 (.Y(n3846), 
	.B(n3455), 
	.A(n4841));
   NAND3X1TS U4097 (.Y(n3756), 
	.C(n3828), 
	.B(\router/data_from_fir ), 
	.A(n3843));
   INVX2TS U4098 (.Y(n4638), 
	.A(n4462));
   INVX2TS U4099 (.Y(n4824), 
	.A(n4648));
   OAI21X1TS U4102 (.Y(n4080), 
	.B0(n4082), 
	.A1(n4078), 
	.A0(n7380));
   OAI21X1TS U4104 (.Y(n4065), 
	.B0(n4067), 
	.A1(n4063), 
	.A0(n7356));
   OAI21X1TS U4108 (.Y(n4130), 
	.B0(n4132), 
	.A1(n7444), 
	.A0(n7450));
   OAI21X1TS U4110 (.Y(n3955), 
	.B0(n3957), 
	.A1(n7335), 
	.A0(n7341));
   OAI21X1TS U4113 (.Y(n3905), 
	.B0(n3907), 
	.A1(n3903), 
	.A0(n7271));
   OAI21X1TS U4114 (.Y(n3890), 
	.B0(n3892), 
	.A1(n3888), 
	.A0(n7247));
   OR2X2TS U4117 (.Y(n4026), 
	.B(\fifo_to_fir/hold[1] ), 
	.A(n5206));
   NOR4XLTS U4118 (.Y(n5206), 
	.D(n5207), 
	.C(\fifo_to_fir/fifo_cell1/controller/valid_read ), 
	.B(\fifo_to_fir/fifo_cell1/controller/write_enable ), 
	.A(n7450));
   OR2X2TS U4119 (.Y(n3851), 
	.B(\fifo_to_fft/hold[1] ), 
	.A(n5248));
   NOR4XLTS U4120 (.Y(n5248), 
	.D(n5249), 
	.C(\fifo_to_fft/fifo_cell1/controller/valid_read ), 
	.B(\fifo_to_fft/fifo_cell1/controller/write_enable ), 
	.A(n7341));
   AOI31X1TS U4122 (.Y(n4032), 
	.B0(\fifo_to_fir/hold[3] ), 
	.A2(n5203), 
	.A1(\fifo_to_fir/fifo_cell3/data_out/N35 ), 
	.A0(n4122));
   NOR3X1TS U4123 (.Y(n4122), 
	.C(n4176), 
	.B(n4175), 
	.A(n8784));
   INVX2TS U4124 (.Y(n4173), 
	.A(n4032));
   NOR3X1TS U4126 (.Y(n3947), 
	.C(n4001), 
	.B(n4000), 
	.A(n8805));
   INVX2TS U4127 (.Y(n3998), 
	.A(n3857));
   AOI31X1TS U4128 (.Y(n4034), 
	.B0(\fifo_to_fir/hold[4] ), 
	.A2(n5202), 
	.A1(\fifo_to_fir/fifo_cell4/data_out/N35 ), 
	.A0(n4117));
   NOR3X1TS U4129 (.Y(n4117), 
	.C(n4173), 
	.B(n4172), 
	.A(n8784));
   AOI31X1TS U4130 (.Y(n3859), 
	.B0(\fifo_to_fft/hold[4] ), 
	.A2(n5244), 
	.A1(\fifo_to_fft/fifo_cell4/data_out/N35 ), 
	.A0(n3942));
   NOR3X1TS U4131 (.Y(n3942), 
	.C(n3998), 
	.B(n3997), 
	.A(n8805));
   AOI31X1TS U4132 (.Y(n3861), 
	.B0(\fifo_to_fft/hold[5] ), 
	.A2(n5243), 
	.A1(\fifo_to_fft/fifo_cell5/data_out/N35 ), 
	.A0(n7315));
   NOR3X1TS U4133 (.Y(n5243), 
	.C(\fifo_to_fft/fifo_cell5/controller/valid_read ), 
	.B(\fifo_to_fft/fifo_cell5/controller/write_enable ), 
	.A(n7311));
   AOI31X1TS U4134 (.Y(n4040), 
	.B0(\fifo_to_fir/hold[7] ), 
	.A2(n5199), 
	.A1(\fifo_to_fir/fifo_cell7/data_out/N35 ), 
	.A0(n4102));
   NOR3X1TS U4135 (.Y(n5199), 
	.C(\fifo_to_fir/fifo_cell7/controller/valid_read ), 
	.B(\fifo_to_fir/fifo_cell7/controller/write_enable ), 
	.A(n7410));
   NOR3X1TS U4136 (.Y(n4102), 
	.C(n4164), 
	.B(n4163), 
	.A(n8785));
   NOR3X1TS U4137 (.Y(n3927), 
	.C(n3989), 
	.B(n3988), 
	.A(n8806));
   AOI31X1TS U4138 (.Y(n4042), 
	.B0(\fifo_to_fir/hold[8] ), 
	.A2(n5198), 
	.A1(\fifo_to_fir/fifo_cell8/data_out/N35 ), 
	.A0(n7404));
   NOR3X1TS U4139 (.Y(n5198), 
	.C(\fifo_to_fir/fifo_cell8/controller/valid_read ), 
	.B(\fifo_to_fir/fifo_cell8/controller/write_enable ), 
	.A(n7400));
   AOI31X1TS U4140 (.Y(n3867), 
	.B0(\fifo_to_fft/hold[8] ), 
	.A2(n5240), 
	.A1(\fifo_to_fft/fifo_cell8/data_out/N35 ), 
	.A0(FE_OFN678_n7295));
   NOR3X1TS U4141 (.Y(n5240), 
	.C(\fifo_to_fft/fifo_cell8/controller/valid_read ), 
	.B(\fifo_to_fft/fifo_cell8/controller/write_enable ), 
	.A(n7291));
   AOI31X1TS U4142 (.Y(n4046), 
	.B0(\fifo_to_fir/hold[10] ), 
	.A2(n5196), 
	.A1(\fifo_to_fir/fifo_cell10/data_out/N35 ), 
	.A0(n4087));
   NOR3X1TS U4143 (.Y(n5196), 
	.C(\fifo_to_fir/fifo_cell10/controller/valid_read ), 
	.B(\fifo_to_fir/fifo_cell10/controller/write_enable ), 
	.A(n7385));
   NOR3X1TS U4144 (.Y(n4087), 
	.C(n4155), 
	.B(n4154), 
	.A(n8786));
   AOI31X1TS U4145 (.Y(n4044), 
	.B0(\fifo_to_fir/hold[9] ), 
	.A2(n5197), 
	.A1(\fifo_to_fir/fifo_cell9/data_out/N35 ), 
	.A0(n7394));
   NOR3X1TS U4146 (.Y(n5197), 
	.C(\fifo_to_fir/fifo_cell9/controller/valid_read ), 
	.B(\fifo_to_fir/fifo_cell9/controller/write_enable ), 
	.A(n7390));
   NOR3X1TS U4147 (.Y(n3912), 
	.C(n3980), 
	.B(n3979), 
	.A(n8807));
   AOI31X1TS U4149 (.Y(n4052), 
	.B0(\fifo_to_fir/hold[13] ), 
	.A2(n5193), 
	.A1(n7365), 
	.A0(\fifo_to_fir/fifo_cell13/data_out/N35 ));
   NOR2BX1TS U4150 (.Y(n3757), 
	.B(n4644), 
	.AN(\router/data_from_iir ));
   NAND2X1TS U4151 (.Y(n4456), 
	.B(n3848), 
	.A(instruction[2]));
   AO21X1TS U4153 (.Y(n3839), 
	.B0(n3838), 
	.A1(n7609), 
	.A0(\router/data_cntl/fir_full_flag ));
   NOR3BX1TS U4165 (.Y(n3720), 
	.C(n3758), 
	.B(n3757), 
	.AN(n3756));
   NAND2X1TS U4192 (.Y(n3458), 
	.B(instruction[31]), 
	.A(instruction[30]));
   OA21XLTS U4193 (.Y(n3794), 
	.B0(n9497), 
	.A1(\fifo_from_fft/fifo_cell0/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell0/controller/f_i_get ));
   OA21XLTS U4194 (.Y(n3774), 
	.B0(n9484), 
	.A1(\fifo_from_fir/fifo_cell0/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell0/controller/f_i_get ));
   NOR3X1TS U4236 (.Y(n4507), 
	.C(n4611), 
	.B(n4610), 
	.A(n8839));
   NOR2X1TS U4241 (.Y(n4508), 
	.B(FE_OFN176_n4507), 
	.A(FE_OFN844_n7619));
   NOR3X1TS U4256 (.Y(n4513), 
	.C(n4614), 
	.B(n4613), 
	.A(n8839));
   NOR3X1TS U4273 (.Y(n4519), 
	.C(n4617), 
	.B(n4616), 
	.A(n8839));
   NOR3X1TS U4284 (.Y(n4525), 
	.C(n4620), 
	.B(n4619), 
	.A(n8838));
   NOR3X1TS U4454 (.Y(n4693), 
	.C(n4797), 
	.B(n4796), 
	.A(n8872));
   NOR2X1TS U4459 (.Y(n4694), 
	.B(FE_OFN518_n4693), 
	.A(FE_OFN846_n7619));
   NOR3X1TS U4474 (.Y(n4699), 
	.C(n4800), 
	.B(n4799), 
	.A(n8872));
   NOR3X1TS U4491 (.Y(n4705), 
	.C(n4803), 
	.B(n4802), 
	.A(n8872));
   NOR3X1TS U4501 (.Y(n4711), 
	.C(n4806), 
	.B(n4805), 
	.A(n8871));
   NOR2X1TS U4520 (.Y(n4718), 
	.B(FE_OFN571_n4717), 
	.A(FE_OFN837_n7619));
   NOR2X1TS U4553 (.Y(n4730), 
	.B(FE_OFN608_n4729), 
	.A(FE_OFN845_n7619));
   NOR3X1TS U4568 (.Y(n4735), 
	.C(n4818), 
	.B(n4817), 
	.A(n8870));
   NOR3X1TS U4583 (.Y(n4741), 
	.C(n4821), 
	.B(n4820), 
	.A(n8870));
   NOR3X1TS U4600 (.Y(n4747), 
	.C(n4824), 
	.B(n4823), 
	.A(n8870));
   NOR2X1TS U4640 (.Y(n3776), 
	.B(n8877), 
	.A(n3772));
   INVX2TS U4643 (.Y(n9433), 
	.A(FE_OFN979_n9462));
   ADDHXLTS U4647 (.S(\router/addr_calc/iir_write_calc/counter/N76 ), 
	.CO(\add_x_22_5/carry[31] ), 
	.B(\add_x_22_5/carry[30] ), 
	.A(\router/addr_calc/iir_write_calc/count[30] ));
   OA21XLTS U4660 (.Y(n4492), 
	.B0(n9483), 
	.A1(\fifo_from_fft/fifo_cell15/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell15/controller/f_i_get ));
   OA21XLTS U4661 (.Y(n4498), 
	.B0(n9483), 
	.A1(\fifo_from_fft/fifo_cell14/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell14/controller/f_i_get ));
   OA21XLTS U4662 (.Y(n4504), 
	.B0(n9483), 
	.A1(\fifo_from_fft/fifo_cell13/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell13/controller/f_i_get ));
   OA21XLTS U4663 (.Y(n4510), 
	.B0(n9483), 
	.A1(\fifo_from_fft/fifo_cell12/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell12/controller/f_i_get ));
   OA21XLTS U4664 (.Y(n4534), 
	.B0(n9482), 
	.A1(\fifo_from_fft/fifo_cell8/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell8/controller/f_i_get ));
   OA21XLTS U4665 (.Y(n4540), 
	.B0(n9481), 
	.A1(\fifo_from_fft/fifo_cell7/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell7/controller/f_i_get ));
   OA21XLTS U4666 (.Y(n4546), 
	.B0(n9481), 
	.A1(\fifo_from_fft/fifo_cell6/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell6/controller/f_i_get ));
   OA21XLTS U4667 (.Y(n4552), 
	.B0(n9481), 
	.A1(\fifo_from_fft/fifo_cell5/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell5/controller/f_i_get ));
   OA21XLTS U4668 (.Y(n4564), 
	.B0(n9481), 
	.A1(\fifo_from_fft/fifo_cell3/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell3/controller/f_i_get ));
   OA21XLTS U4669 (.Y(n4570), 
	.B0(n9497), 
	.A1(\fifo_from_fft/fifo_cell2/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell2/controller/f_i_get ));
   NAND2X1TS U4670 (.Y(n4572), 
	.B(\fifo_from_fft/fifo_cell1/reg_gtok/token ), 
	.A(FE_OFN721_n4643));
   NAND2X1TS U4671 (.Y(n4566), 
	.B(\fifo_from_fft/fifo_cell2/reg_gtok/token ), 
	.A(FE_OFN719_n4643));
   NAND2X1TS U4672 (.Y(n4560), 
	.B(\fifo_from_fft/fifo_cell3/reg_gtok/token ), 
	.A(n4643));
   NAND2X1TS U4673 (.Y(n4554), 
	.B(\fifo_from_fft/fifo_cell4/reg_gtok/token ), 
	.A(FE_OFN1823_n4643));
   NAND2X1TS U4674 (.Y(n4548), 
	.B(\fifo_from_fft/fifo_cell5/reg_gtok/token ), 
	.A(FE_OFN720_n4643));
   NAND2X1TS U4675 (.Y(n4542), 
	.B(\fifo_from_fft/fifo_cell6/reg_gtok/token ), 
	.A(FE_OFN723_n4643));
   NAND2X1TS U4676 (.Y(n4536), 
	.B(\fifo_from_fft/fifo_cell7/reg_gtok/token ), 
	.A(FE_OFN727_n4643));
   NAND2X1TS U4677 (.Y(n4530), 
	.B(\fifo_from_fft/fifo_cell8/reg_gtok/token ), 
	.A(FE_OFN727_n4643));
   NAND2X1TS U4678 (.Y(n4524), 
	.B(\fifo_from_fft/fifo_cell9/reg_gtok/token ), 
	.A(FE_OFN726_n4643));
   NAND2X1TS U4679 (.Y(n4518), 
	.B(\fifo_from_fft/fifo_cell10/reg_gtok/token ), 
	.A(FE_OFN726_n4643));
   NAND2X1TS U4680 (.Y(n4512), 
	.B(\fifo_from_fft/fifo_cell11/reg_gtok/token ), 
	.A(FE_OFN728_n4643));
   OA21XLTS U4681 (.Y(n4131), 
	.B0(n9492), 
	.A1(\fifo_to_fir/fifo_cell1/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell1/controller/f_i_get ));
   NAND2X1TS U4682 (.Y(n4123), 
	.B(n4134), 
	.A(\fifo_to_fir/fifo_cell1/reg_gtok/token ));
   OA21XLTS U4683 (.Y(n4126), 
	.B0(n9492), 
	.A1(\fifo_to_fir/fifo_cell2/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell2/controller/f_i_get ));
   NAND2X1TS U4684 (.Y(n4118), 
	.B(FE_OFN686_n4134), 
	.A(\fifo_to_fir/fifo_cell2/reg_gtok/token ));
   OA21XLTS U4685 (.Y(n4121), 
	.B0(n9493), 
	.A1(\fifo_to_fir/fifo_cell3/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell3/controller/f_i_get ));
   OA21XLTS U4686 (.Y(n4116), 
	.B0(n9493), 
	.A1(\fifo_to_fir/fifo_cell4/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell4/controller/f_i_get ));
   NAND2X1TS U4687 (.Y(n4108), 
	.B(FE_OFN687_n4134), 
	.A(\fifo_to_fir/fifo_cell4/reg_gtok/token ));
   OA21XLTS U4688 (.Y(n4111), 
	.B0(n9493), 
	.A1(\fifo_to_fir/fifo_cell5/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell5/controller/f_i_get ));
   NAND2X1TS U4689 (.Y(n4103), 
	.B(FE_OFN687_n4134), 
	.A(\fifo_to_fir/fifo_cell5/reg_gtok/token ));
   OA21XLTS U4690 (.Y(n4106), 
	.B0(n9493), 
	.A1(\fifo_to_fir/fifo_cell6/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell6/controller/f_i_get ));
   NAND2X1TS U4691 (.Y(n4098), 
	.B(FE_OFN688_n4134), 
	.A(\fifo_to_fir/fifo_cell6/reg_gtok/token ));
   OA21XLTS U4692 (.Y(n4101), 
	.B0(n9494), 
	.A1(\fifo_to_fir/fifo_cell7/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell7/controller/f_i_get ));
   NAND2X1TS U4693 (.Y(n4093), 
	.B(FE_OFN688_n4134), 
	.A(\fifo_to_fir/fifo_cell7/reg_gtok/token ));
   OA21XLTS U4694 (.Y(n4096), 
	.B0(n9494), 
	.A1(\fifo_to_fir/fifo_cell8/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell8/controller/f_i_get ));
   NAND2X1TS U4695 (.Y(n4088), 
	.B(FE_OFN689_n4134), 
	.A(\fifo_to_fir/fifo_cell8/reg_gtok/token ));
   OA21XLTS U4696 (.Y(n4091), 
	.B0(n9494), 
	.A1(\fifo_to_fir/fifo_cell9/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell9/controller/f_i_get ));
   NAND2X1TS U4697 (.Y(n4083), 
	.B(FE_OFN692_n4134), 
	.A(\fifo_to_fir/fifo_cell9/reg_gtok/token ));
   OA21XLTS U4698 (.Y(n4086), 
	.B0(n9494), 
	.A1(\fifo_to_fir/fifo_cell10/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell10/controller/f_i_get ));
   NAND2X1TS U4699 (.Y(n4078), 
	.B(FE_OFN694_n4134), 
	.A(\fifo_to_fir/fifo_cell10/reg_gtok/token ));
   OA21XLTS U4700 (.Y(n4081), 
	.B0(n9495), 
	.A1(\fifo_to_fir/fifo_cell11/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell11/controller/f_i_get ));
   NAND2X1TS U4701 (.Y(n4073), 
	.B(FE_OFN694_n4134), 
	.A(\fifo_to_fir/fifo_cell11/reg_gtok/token ));
   OA21XLTS U4702 (.Y(n4076), 
	.B0(n9495), 
	.A1(\fifo_to_fir/fifo_cell12/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell12/controller/f_i_get ));
   NAND2X1TS U4703 (.Y(n4068), 
	.B(FE_OFN695_n4134), 
	.A(\fifo_to_fir/fifo_cell12/reg_gtok/token ));
   OA21XLTS U4704 (.Y(n4071), 
	.B0(n9495), 
	.A1(\fifo_to_fir/fifo_cell13/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell13/controller/f_i_get ));
   NAND2X1TS U4705 (.Y(n4063), 
	.B(FE_OFN695_n4134), 
	.A(\fifo_to_fir/fifo_cell13/reg_gtok/token ));
   OA21XLTS U4706 (.Y(n4066), 
	.B0(n9495), 
	.A1(\fifo_to_fir/fifo_cell14/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell14/controller/f_i_get ));
   OA21XLTS U4707 (.Y(n4061), 
	.B0(n9496), 
	.A1(\fifo_to_fir/fifo_cell15/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell15/controller/f_i_get ));
   OA21XLTS U4708 (.Y(n3809), 
	.B0(n9492), 
	.A1(\fifo_to_fir/fifo_cell0/controller/f_i_put ), 
	.A0(\fifo_to_fir/fifo_cell0/controller/f_i_get ));
   OA21XLTS U4710 (.Y(n3956), 
	.B0(n9488), 
	.A1(\fifo_to_fft/fifo_cell1/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell1/controller/f_i_get ));
   NAND2X1TS U4711 (.Y(n3948), 
	.B(FE_OFN701_n3959), 
	.A(\fifo_to_fft/fifo_cell1/reg_gtok/token ));
   OA21XLTS U4712 (.Y(n3951), 
	.B0(n9488), 
	.A1(\fifo_to_fft/fifo_cell2/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell2/controller/f_i_get ));
   NAND2X1TS U4713 (.Y(n3943), 
	.B(FE_OFN704_n3959), 
	.A(\fifo_to_fft/fifo_cell2/reg_gtok/token ));
   OA21XLTS U4714 (.Y(n3946), 
	.B0(n9489), 
	.A1(\fifo_to_fft/fifo_cell3/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell3/controller/f_i_get ));
   NAND2X1TS U4715 (.Y(n3938), 
	.B(FE_OFN704_n3959), 
	.A(\fifo_to_fft/fifo_cell3/reg_gtok/token ));
   OA21XLTS U4716 (.Y(n3941), 
	.B0(n9489), 
	.A1(\fifo_to_fft/fifo_cell4/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell4/controller/f_i_get ));
   NAND2X1TS U4717 (.Y(n3933), 
	.B(FE_OFN708_n3959), 
	.A(\fifo_to_fft/fifo_cell4/reg_gtok/token ));
   OA21XLTS U4718 (.Y(n3936), 
	.B0(n9489), 
	.A1(\fifo_to_fft/fifo_cell5/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell5/controller/f_i_get ));
   NAND2X1TS U4719 (.Y(n3928), 
	.B(FE_OFN705_n3959), 
	.A(\fifo_to_fft/fifo_cell5/reg_gtok/token ));
   OA21XLTS U4720 (.Y(n3931), 
	.B0(n9496), 
	.A1(\fifo_to_fft/fifo_cell6/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell6/controller/f_i_get ));
   NAND2X1TS U4721 (.Y(n3923), 
	.B(FE_OFN705_n3959), 
	.A(\fifo_to_fft/fifo_cell6/reg_gtok/token ));
   OA21XLTS U4722 (.Y(n3926), 
	.B0(n9490), 
	.A1(\fifo_to_fft/fifo_cell7/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell7/controller/f_i_get ));
   NAND2X1TS U4723 (.Y(n3918), 
	.B(FE_OFN702_n3959), 
	.A(\fifo_to_fft/fifo_cell7/reg_gtok/token ));
   OA21XLTS U4724 (.Y(n3921), 
	.B0(n9490), 
	.A1(\fifo_to_fft/fifo_cell8/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell8/controller/f_i_get ));
   NAND2X1TS U4726 (.Y(n3913), 
	.B(FE_OFN702_n3959), 
	.A(\fifo_to_fft/fifo_cell8/reg_gtok/token ));
   OA21XLTS U4727 (.Y(n3916), 
	.B0(n9490), 
	.A1(\fifo_to_fft/fifo_cell9/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell9/controller/f_i_get ));
   NAND2X1TS U4728 (.Y(n3908), 
	.B(FE_OFN706_n3959), 
	.A(\fifo_to_fft/fifo_cell9/reg_gtok/token ));
   OA21XLTS U4729 (.Y(n3911), 
	.B0(n9490), 
	.A1(\fifo_to_fft/fifo_cell10/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell10/controller/f_i_get ));
   NAND2X1TS U4730 (.Y(n3903), 
	.B(FE_OFN707_n3959), 
	.A(\fifo_to_fft/fifo_cell10/reg_gtok/token ));
   OA21XLTS U4731 (.Y(n3906), 
	.B0(n9491), 
	.A1(\fifo_to_fft/fifo_cell11/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell11/controller/f_i_get ));
   NAND2X1TS U4732 (.Y(n3898), 
	.B(FE_OFN707_n3959), 
	.A(\fifo_to_fft/fifo_cell11/reg_gtok/token ));
   OA21XLTS U4733 (.Y(n3901), 
	.B0(n9491), 
	.A1(\fifo_to_fft/fifo_cell12/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell12/controller/f_i_get ));
   NAND2X1TS U4734 (.Y(n3893), 
	.B(FE_OFN703_n3959), 
	.A(\fifo_to_fft/fifo_cell12/reg_gtok/token ));
   OA21XLTS U4735 (.Y(n3896), 
	.B0(n9491), 
	.A1(\fifo_to_fft/fifo_cell13/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell13/controller/f_i_get ));
   NAND2X1TS U4736 (.Y(n3888), 
	.B(FE_OFN699_n3959), 
	.A(\fifo_to_fft/fifo_cell13/reg_gtok/token ));
   OA21XLTS U4737 (.Y(n3891), 
	.B0(n9491), 
	.A1(\fifo_to_fft/fifo_cell14/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell14/controller/f_i_get ));
   OA21XLTS U4738 (.Y(n3886), 
	.B0(n9492), 
	.A1(\fifo_to_fft/fifo_cell15/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell15/controller/f_i_get ));
   OA21XLTS U4739 (.Y(n3820), 
	.B0(n9488), 
	.A1(\fifo_to_fft/fifo_cell0/controller/f_i_put ), 
	.A0(\fifo_to_fft/fifo_cell0/controller/f_i_get ));
   OA21XLTS U4748 (.Y(n4678), 
	.B0(n9487), 
	.A1(\fifo_from_fir/fifo_cell15/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell15/controller/f_i_get ));
   OA21XLTS U4749 (.Y(n4720), 
	.B0(n9486), 
	.A1(\fifo_from_fir/fifo_cell8/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell8/controller/f_i_get ));
   OA21XLTS U4750 (.Y(n4726), 
	.B0(n9485), 
	.A1(\fifo_from_fir/fifo_cell7/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell7/controller/f_i_get ));
   OA21XLTS U4751 (.Y(n4732), 
	.B0(n9485), 
	.A1(\fifo_from_fir/fifo_cell6/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell6/controller/f_i_get ));
   OA21XLTS U4752 (.Y(n4738), 
	.B0(n9485), 
	.A1(\fifo_from_fir/fifo_cell5/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell5/controller/f_i_get ));
   OA21XLTS U4753 (.Y(n4744), 
	.B0(n9485), 
	.A1(\fifo_from_fir/fifo_cell4/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell4/controller/f_i_get ));
   NAND2X1TS U4754 (.Y(n4758), 
	.B(\fifo_from_fir/fifo_cell1/reg_gtok/token ), 
	.A(n4829));
   NAND2X1TS U4755 (.Y(n4752), 
	.B(\fifo_from_fir/fifo_cell2/reg_gtok/token ), 
	.A(FE_OFN737_n4829));
   NAND2X1TS U4756 (.Y(n4746), 
	.B(\fifo_from_fir/fifo_cell3/reg_gtok/token ), 
	.A(FE_OFN738_n4829));
   NAND2X1TS U4757 (.Y(n4740), 
	.B(\fifo_from_fir/fifo_cell4/reg_gtok/token ), 
	.A(FE_OFN740_n4829));
   NAND2X1TS U4758 (.Y(n4734), 
	.B(\fifo_from_fir/fifo_cell5/reg_gtok/token ), 
	.A(FE_OFN743_n4829));
   NAND2X1TS U4759 (.Y(n4728), 
	.B(\fifo_from_fir/fifo_cell6/reg_gtok/token ), 
	.A(FE_OFN743_n4829));
   NAND2X1TS U4760 (.Y(n4722), 
	.B(\fifo_from_fir/fifo_cell7/reg_gtok/token ), 
	.A(FE_OFN744_n4829));
   NAND2X1TS U4761 (.Y(n4716), 
	.B(\fifo_from_fir/fifo_cell8/reg_gtok/token ), 
	.A(FE_OFN744_n4829));
   NAND2X1TS U4762 (.Y(n4710), 
	.B(\fifo_from_fir/fifo_cell9/reg_gtok/token ), 
	.A(FE_OFN739_n4829));
   NAND2X1TS U4763 (.Y(n4704), 
	.B(\fifo_from_fir/fifo_cell10/reg_gtok/token ), 
	.A(FE_OFN739_n4829));
   NAND2X1TS U4764 (.Y(n4698), 
	.B(\fifo_from_fir/fifo_cell11/reg_gtok/token ), 
	.A(FE_OFN741_n4829));
   INVX2TS U4810 (.Y(n8838), 
	.A(FE_OFN697_n8052));
   INVX2TS U4811 (.Y(n8871), 
	.A(FE_OFN679_n8050));
   NOR3X1TS U4816 (.Y(n4561), 
	.C(n4638), 
	.B(n4637), 
	.A(n8837));
   INVX2TS U4831 (.Y(n9465), 
	.A(FE_OFN833_n7619));
   NAND2X1TS U4832 (.Y(n3486), 
	.B(\router/addr_calc/iir_write_calc/counter/N40 ), 
	.A(\router/data_from_iir ));
   INVX2TS U4833 (.Y(n9480), 
	.A(FE_OFN782_n7619));
   INVX2TS U4835 (.Y(n9497), 
	.A(FE_OFN813_n7619));
   INVX2TS U4836 (.Y(n9406), 
	.A(FE_OFN988_n9431));
   INVX2TS U4837 (.Y(n9432), 
	.A(FE_OFN976_n9462));
   INVX2TS U4838 (.Y(n9407), 
	.A(FE_OFN986_n9431));
   INVX2TS U4839 (.Y(n9514), 
	.A(FE_OFN789_n7619));
   INVX2TS U4840 (.Y(n9435), 
	.A(n9462));
   INVX2TS U4841 (.Y(n8376), 
	.A(n8055));
   INVX2TS U4842 (.Y(n8711), 
	.A(n8054));
   INVX2TS U4847 (.Y(n8472), 
	.A(n8056));
   INVX2TS U4849 (.Y(n8137), 
	.A(FE_OFN664_n8053));
   AND2X2TS U4876 (.Y(n5702), 
	.B(FE_OFN715_n4207), 
	.A(\mips/mips/accbypass ));
   AND2X2TS U4877 (.Y(n5584), 
	.B(\mips/mips/accfullinstruction[21] ), 
	.A(FE_OFN713_n4207));
   AND2X2TS U4878 (.Y(n5585), 
	.B(\mips/mips/accfullinstruction[20] ), 
	.A(FE_OFN713_n4207));
   AND2X2TS U4879 (.Y(n5586), 
	.B(\mips/mips/accfullinstruction[19] ), 
	.A(FE_OFN716_n4207));
   AND2X2TS U4880 (.Y(n5587), 
	.B(\mips/mips/accfullinstruction[18] ), 
	.A(FE_OFN716_n4207));
   AND2X2TS U4881 (.Y(n5588), 
	.B(\mips/mips/accfullinstruction[17] ), 
	.A(FE_OFN716_n4207));
   AND2X2TS U4882 (.Y(n5589), 
	.B(\mips/mips/accfullinstruction[16] ), 
	.A(FE_OFN713_n4207));
   AND2X2TS U4883 (.Y(n5590), 
	.B(\mips/mips/accfullinstruction[15] ), 
	.A(FE_OFN714_n4207));
   AND2X2TS U4884 (.Y(n5591), 
	.B(\mips/mips/accfullinstruction[14] ), 
	.A(FE_OFN716_n4207));
   AND2X2TS U4885 (.Y(n5592), 
	.B(\mips/mips/accfullinstruction[13] ), 
	.A(FE_OFN712_n4207));
   AND2X2TS U4886 (.Y(n5593), 
	.B(\mips/mips/accfullinstruction[12] ), 
	.A(FE_OFN715_n4207));
   AND2X2TS U4887 (.Y(n5594), 
	.B(\mips/mips/accfullinstruction[11] ), 
	.A(FE_OFN714_n4207));
   AND2X2TS U4888 (.Y(n5595), 
	.B(\mips/mips/accfullinstruction[10] ), 
	.A(FE_OFN715_n4207));
   AND2X2TS U4889 (.Y(n5596), 
	.B(\mips/mips/accfullinstruction[9] ), 
	.A(FE_OFN712_n4207));
   AND2X2TS U4890 (.Y(n5597), 
	.B(\mips/mips/accfullinstruction[8] ), 
	.A(FE_OFN709_n4207));
   AND2X2TS U4891 (.Y(n5598), 
	.B(\mips/mips/accfullinstruction[7] ), 
	.A(FE_OFN710_n4207));
   AND2X2TS U4892 (.Y(n5599), 
	.B(\mips/mips/accfullinstruction[6] ), 
	.A(FE_OFN711_n4207));
   AND2X2TS U4893 (.Y(n5601), 
	.B(\mips/mips/accfullinstruction[4] ), 
	.A(n4207));
   AND2X2TS U4894 (.Y(n5604), 
	.B(\mips/mips/accfullinstruction[1] ), 
	.A(n4207));
   AND2X2TS U4895 (.Y(n5605), 
	.B(\mips/mips/accfullinstruction[0] ), 
	.A(FE_OFN715_n4207));
   AOI222XLTS U5208 (.Y(n3751), 
	.C1(fir_data_in[2]), 
	.C0(FE_OFN747_n3722), 
	.B1(FE_MDBN5_), 
	.B0(FE_OFN757_n3721), 
	.A1(\router/data_cntl/data_in[2] ), 
	.A0(FE_OFN768_n3720));
   AOI222XLTS U5209 (.Y(n3750), 
	.C1(fir_data_in[3]), 
	.C0(FE_OFN750_n3722), 
	.B1(FE_MDBN6_), 
	.B0(FE_OFN760_n3721), 
	.A1(\router/data_cntl/data_in[3] ), 
	.A0(FE_OFN771_n3720));
   AOI222XLTS U5210 (.Y(n3748), 
	.C1(fir_data_in[5]), 
	.C0(FE_OFN749_n3722), 
	.B1(FE_MDBN7_), 
	.B0(FE_OFN759_n3721), 
	.A1(\router/data_cntl/data_in[5] ), 
	.A0(FE_OFN770_n3720));
   AOI222XLTS U5211 (.Y(n3747), 
	.C1(fir_data_in[6]), 
	.C0(FE_OFN747_n3722), 
	.B1(fft_data_in[6]), 
	.B0(FE_OFN757_n3721), 
	.A1(\router/data_cntl/data_in[6] ), 
	.A0(FE_OFN768_n3720));
   AOI222XLTS U5212 (.Y(n3745), 
	.C1(fir_data_in[8]), 
	.C0(FE_OFN754_n3722), 
	.B1(fft_data_in[8]), 
	.B0(FE_OFN764_n3721), 
	.A1(\router/data_cntl/data_in[8] ), 
	.A0(FE_OFN775_n3720));
   AOI222XLTS U5213 (.Y(n3744), 
	.C1(fir_data_in[9]), 
	.C0(FE_OFN754_n3722), 
	.B1(fft_data_in[9]), 
	.B0(FE_OFN764_n3721), 
	.A1(\router/data_cntl/data_in[9] ), 
	.A0(FE_OFN775_n3720));
   AOI222XLTS U5214 (.Y(n3741), 
	.C1(fir_data_in[12]), 
	.C0(FE_OFN750_n3722), 
	.B1(fft_data_in[12]), 
	.B0(FE_OFN760_n3721), 
	.A1(\router/data_cntl/data_in[12] ), 
	.A0(FE_OFN771_n3720));
   AOI222XLTS U5215 (.Y(n3740), 
	.C1(fir_data_in[13]), 
	.C0(FE_OFN753_n3722), 
	.B1(fft_data_in[13]), 
	.B0(FE_OFN763_n3721), 
	.A1(\router/data_cntl/data_in[13] ), 
	.A0(FE_OFN774_n3720));
   AOI222XLTS U5216 (.Y(n3739), 
	.C1(fir_data_in[14]), 
	.C0(FE_OFN751_n3722), 
	.B1(fft_data_in[14]), 
	.B0(FE_OFN761_n3721), 
	.A1(\router/data_cntl/data_in[14] ), 
	.A0(FE_OFN772_n3720));
   AOI222XLTS U5217 (.Y(n3738), 
	.C1(fir_data_in[15]), 
	.C0(FE_OFN753_n3722), 
	.B1(fft_data_in[15]), 
	.B0(FE_OFN763_n3721), 
	.A1(\router/data_cntl/data_in[15] ), 
	.A0(FE_OFN774_n3720));
   AOI222XLTS U5218 (.Y(n3737), 
	.C1(fir_data_in[16]), 
	.C0(FE_OFN746_n3722), 
	.B1(fft_data_in[16]), 
	.B0(FE_OFN755_n3721), 
	.A1(\router/data_cntl/data_in[16] ), 
	.A0(FE_OFN767_n3720));
   AOI222XLTS U5219 (.Y(n3736), 
	.C1(fir_data_in[17]), 
	.C0(FE_OFN746_n3722), 
	.B1(fft_data_in[17]), 
	.B0(FE_OFN755_n3721), 
	.A1(\router/data_cntl/data_in[17] ), 
	.A0(FE_OFN767_n3720));
   AOI222XLTS U5220 (.Y(n3735), 
	.C1(fir_data_in[18]), 
	.C0(FE_OFN753_n3722), 
	.B1(fft_data_in[18]), 
	.B0(FE_OFN763_n3721), 
	.A1(\router/data_cntl/data_in[18] ), 
	.A0(FE_OFN774_n3720));
   AOI222XLTS U5221 (.Y(n3729), 
	.C1(fir_data_in[24]), 
	.C0(FE_OFN749_n3722), 
	.B1(FE_MDBN8_), 
	.B0(FE_OFN759_n3721), 
	.A1(\router/data_cntl/data_in[24] ), 
	.A0(FE_OFN770_n3720));
   AOI222XLTS U5222 (.Y(n3728), 
	.C1(fir_data_in[25]), 
	.C0(FE_OFN749_n3722), 
	.B1(fft_data_in[25]), 
	.B0(FE_OFN759_n3721), 
	.A1(\router/data_cntl/data_in[25] ), 
	.A0(FE_OFN770_n3720));
   AOI222XLTS U5223 (.Y(n3727), 
	.C1(fir_data_in[26]), 
	.C0(FE_OFN748_n3722), 
	.B1(FE_MDBN9_), 
	.B0(FE_OFN758_n3721), 
	.A1(\router/data_cntl/data_in[26] ), 
	.A0(FE_OFN769_n3720));
   NAND2X1TS U5228 (.Y(n5250), 
	.B(\fifo_to_fft/tok_xnor_put ), 
	.A(\fifo_to_fft/fifo_cell0/reg_ptok/N29 ));
   NAND2X1TS U5229 (.Y(n5208), 
	.B(\fifo_to_fir/tok_xnor_put ), 
	.A(\fifo_to_fir/fifo_cell0/reg_ptok/N29 ));
   NAND2X1TS U5230 (.Y(n5327), 
	.B(\fifo_from_fft/tok_xnor_put ), 
	.A(\fifo_from_fft/fifo_cell0/reg_ptok/N29 ));
   INVX2TS U5231 (.Y(n8844), 
	.A(n8052));
   NAND2X1TS U5232 (.Y(n5288), 
	.B(\fifo_from_fir/tok_xnor_put ), 
	.A(\fifo_from_fir/fifo_cell0/reg_ptok/N29 ));
   INVX2TS U5233 (.Y(n8877), 
	.A(FE_OFN681_n8050));
   NOR2X1TS U5234 (.Y(n3957), 
	.B(n5250), 
	.A(n8812));
   INVX2TS U5235 (.Y(\fifo_to_fft/fifo_cell1/data_out/N35 ), 
	.A(n7335));
   NOR2X1TS U5236 (.Y(n4132), 
	.B(n5208), 
	.A(n8791));
   INVX2TS U5237 (.Y(\fifo_to_fir/fifo_cell1/data_out/N35 ), 
	.A(n7444));
   INVX2TS U5241 (.Y(\fifo_from_fft/fifo_cell2/data_out/N35 ), 
	.A(n4572));
   INVX2TS U5242 (.Y(\fifo_from_fft/fifo_cell3/data_out/N35 ), 
	.A(n4566));
   INVX2TS U5243 (.Y(\fifo_from_fft/fifo_cell4/data_out/N35 ), 
	.A(n4560));
   INVX2TS U5244 (.Y(\fifo_from_fft/fifo_cell5/data_out/N35 ), 
	.A(n4554));
   INVX2TS U5245 (.Y(\fifo_from_fft/fifo_cell6/data_out/N35 ), 
	.A(n4548));
   INVX2TS U5246 (.Y(\fifo_from_fft/fifo_cell7/data_out/N35 ), 
	.A(n4542));
   INVX2TS U5247 (.Y(\fifo_from_fft/fifo_cell8/data_out/N35 ), 
	.A(n4536));
   INVX2TS U5248 (.Y(\fifo_from_fft/fifo_cell9/data_out/N35 ), 
	.A(n4530));
   INVX2TS U5249 (.Y(\fifo_from_fft/fifo_cell10/data_out/N35 ), 
	.A(n4524));
   INVX2TS U5250 (.Y(\fifo_from_fft/fifo_cell11/data_out/N35 ), 
	.A(n4518));
   INVX2TS U5251 (.Y(\fifo_from_fft/fifo_cell12/data_out/N35 ), 
	.A(n4512));
   INVX2TS U5252 (.Y(\fifo_to_fir/fifo_cell3/data_out/N35 ), 
	.A(n4118));
   INVX2TS U5253 (.Y(\fifo_to_fir/fifo_cell5/data_out/N35 ), 
	.A(n4108));
   INVX2TS U5254 (.Y(\fifo_to_fir/fifo_cell6/data_out/N35 ), 
	.A(n4103));
   INVX2TS U5255 (.Y(\fifo_to_fir/fifo_cell7/data_out/N35 ), 
	.A(n4098));
   INVX2TS U5256 (.Y(\fifo_to_fir/fifo_cell8/data_out/N35 ), 
	.A(n4093));
   INVX2TS U5257 (.Y(\fifo_to_fir/fifo_cell9/data_out/N35 ), 
	.A(n4088));
   INVX2TS U5258 (.Y(\fifo_to_fir/fifo_cell10/data_out/N35 ), 
	.A(n4083));
   INVX2TS U5259 (.Y(\fifo_to_fir/fifo_cell11/data_out/N35 ), 
	.A(n4078));
   INVX2TS U5260 (.Y(\fifo_to_fir/fifo_cell12/data_out/N35 ), 
	.A(n4073));
   INVX2TS U5261 (.Y(\fifo_to_fir/fifo_cell13/data_out/N35 ), 
	.A(n4068));
   INVX2TS U5263 (.Y(\fifo_to_fir/fifo_cell14/data_out/N35 ), 
	.A(n4063));
   AO21X1TS U5264 (.Y(n8095), 
	.B0(n3825), 
	.A1(n3474), 
	.A0(n3826));
   INVX2TS U5265 (.Y(\fifo_to_fft/fifo_cell3/data_out/N35 ), 
	.A(n3943));
   INVX2TS U5266 (.Y(\fifo_to_fft/fifo_cell4/data_out/N35 ), 
	.A(n3938));
   INVX2TS U5267 (.Y(\fifo_to_fft/fifo_cell5/data_out/N35 ), 
	.A(n3933));
   INVX2TS U5268 (.Y(\fifo_to_fft/fifo_cell6/data_out/N35 ), 
	.A(n3928));
   INVX2TS U5269 (.Y(\fifo_to_fft/fifo_cell7/data_out/N35 ), 
	.A(n3923));
   INVX2TS U5270 (.Y(\fifo_to_fft/fifo_cell8/data_out/N35 ), 
	.A(n3918));
   INVX2TS U5271 (.Y(\fifo_to_fft/fifo_cell9/data_out/N35 ), 
	.A(n3913));
   INVX2TS U5272 (.Y(\fifo_to_fft/fifo_cell10/data_out/N35 ), 
	.A(n3908));
   INVX2TS U5273 (.Y(\fifo_to_fft/fifo_cell11/data_out/N35 ), 
	.A(n3903));
   INVX2TS U5274 (.Y(\fifo_to_fft/fifo_cell12/data_out/N35 ), 
	.A(n3898));
   INVX2TS U5275 (.Y(\fifo_to_fft/fifo_cell13/data_out/N35 ), 
	.A(n3893));
   INVX2TS U5277 (.Y(\fifo_to_fft/fifo_cell14/data_out/N35 ), 
	.A(n3888));
   INVX2TS U5282 (.Y(\fifo_from_fir/fifo_cell2/data_out/N35 ), 
	.A(n4758));
   INVX2TS U5283 (.Y(\fifo_from_fir/fifo_cell3/data_out/N35 ), 
	.A(n4752));
   INVX2TS U5284 (.Y(\fifo_from_fir/fifo_cell4/data_out/N35 ), 
	.A(n4746));
   INVX2TS U5285 (.Y(\fifo_from_fir/fifo_cell5/data_out/N35 ), 
	.A(n4740));
   INVX2TS U5286 (.Y(\fifo_from_fir/fifo_cell6/data_out/N35 ), 
	.A(n4734));
   INVX2TS U5287 (.Y(\fifo_from_fir/fifo_cell7/data_out/N35 ), 
	.A(n4728));
   INVX2TS U5288 (.Y(\fifo_from_fir/fifo_cell8/data_out/N35 ), 
	.A(n4722));
   INVX2TS U5289 (.Y(\fifo_from_fir/fifo_cell9/data_out/N35 ), 
	.A(n4716));
   INVX2TS U5290 (.Y(\fifo_from_fir/fifo_cell10/data_out/N35 ), 
	.A(n4710));
   INVX2TS U5291 (.Y(\fifo_from_fir/fifo_cell11/data_out/N35 ), 
	.A(n4704));
   INVX2TS U5292 (.Y(\fifo_from_fir/fifo_cell12/data_out/N35 ), 
	.A(n4698));
   NOR2X1TS U5294 (.Y(n3777), 
	.B(FE_OFN419_n3776), 
	.A(FE_OFN841_n7619));
   NOR2X1TS U5295 (.Y(n3797), 
	.B(FE_OFN73_n3796), 
	.A(FE_OFN844_n7619));
   NOR2X1TS U5297 (.Y(n3796), 
	.B(n8844), 
	.A(n3792));
   AOI21X1TS U5298 (.Y(n3792), 
	.B0(n3784), 
	.A1(n4488), 
	.A0(\fifo_from_fft/hang[14] ));
   NOR2X1TS U5299 (.Y(n4490), 
	.B(FE_OFN142_n4489), 
	.A(FE_OFN847_n7619));
   AOI31X1TS U5300 (.Y(n4488), 
	.B0(\fifo_from_fft/hold[15] ), 
	.A2(n5312), 
	.A1(n4489), 
	.A0(\fifo_from_fft/fifo_cell15/data_out/N35 ));
   NOR2X1TS U5301 (.Y(n4676), 
	.B(FE_OFN480_n4675), 
	.A(FE_OFN831_n7619));
   NOR3X1TS U5302 (.Y(n4489), 
	.C(n4602), 
	.B(n4601), 
	.A(n8840));
   NOR3X1TS U5305 (.Y(n4675), 
	.C(n4788), 
	.B(n4787), 
	.A(n8873));
   AOI31X1TS U5306 (.Y(n4486), 
	.B0(\fifo_from_fft/hold[14] ), 
	.A2(n5313), 
	.A1(n4495), 
	.A0(\fifo_from_fft/fifo_cell14/data_out/N35 ));
   NOR2X1TS U5307 (.Y(n4496), 
	.B(FE_OFN162_n4495), 
	.A(FE_OFN836_n7619));
   AOI31X1TS U5308 (.Y(n4672), 
	.B0(\fifo_from_fir/hold[14] ), 
	.A2(n5274), 
	.A1(FE_OFN496_n4681), 
	.A0(\fifo_from_fir/fifo_cell14/data_out/N35 ));
   NOR2X1TS U5309 (.Y(n4682), 
	.B(FE_OFN502_n4681), 
	.A(FE_OFN841_n7619));
   NOR3X1TS U5311 (.Y(n4495), 
	.C(n4605), 
	.B(n4604), 
	.A(n8840));
   NOR3X1TS U5313 (.Y(n4681), 
	.C(n4791), 
	.B(n4790), 
	.A(n8873));
   AOI31X1TS U5314 (.Y(n4484), 
	.B0(\fifo_from_fft/hold[13] ), 
	.A2(n5314), 
	.A1(n8711), 
	.A0(\fifo_from_fft/fifo_cell13/data_out/N35 ));
   AOI31X1TS U5315 (.Y(n4670), 
	.B0(\fifo_from_fir/hold[13] ), 
	.A2(n5275), 
	.A1(n8376), 
	.A0(\fifo_from_fir/fifo_cell13/data_out/N35 ));
   AOI31X1TS U5318 (.Y(n4482), 
	.B0(\fifo_from_fft/hold[12] ), 
	.A2(n5315), 
	.A1(\fifo_from_fft/fifo_cell12/data_out/N35 ), 
	.A0(FE_OFN175_n4507));
   AOI31X1TS U5319 (.Y(n4668), 
	.B0(\fifo_from_fir/hold[12] ), 
	.A2(n5276), 
	.A1(\fifo_from_fir/fifo_cell12/data_out/N35 ), 
	.A0(n4693));
   AOI31X1TS U5320 (.Y(n4480), 
	.B0(\fifo_from_fft/hold[11] ), 
	.A2(n5316), 
	.A1(\fifo_from_fft/fifo_cell11/data_out/N35 ), 
	.A0(FE_OFN199_n4513));
   NOR2X1TS U5321 (.Y(n4514), 
	.B(FE_OFN199_n4513), 
	.A(FE_OFN836_n7619));
   AOI31X1TS U5322 (.Y(n4666), 
	.B0(\fifo_from_fir/hold[11] ), 
	.A2(n5277), 
	.A1(\fifo_from_fir/fifo_cell11/data_out/N35 ), 
	.A0(FE_OFN534_n4699));
   NOR2X1TS U5323 (.Y(n4700), 
	.B(n4699), 
	.A(FE_OFN831_n7619));
   AOI31X1TS U5326 (.Y(n4478), 
	.B0(\fifo_from_fft/hold[10] ), 
	.A2(n5317), 
	.A1(\fifo_from_fft/fifo_cell10/data_out/N35 ), 
	.A0(FE_OFN209_n4519));
   NOR2X1TS U5327 (.Y(n4706), 
	.B(FE_OFN547_n4705), 
	.A(FE_OFN846_n7619));
   AOI31X1TS U5328 (.Y(n4664), 
	.B0(\fifo_from_fir/hold[10] ), 
	.A2(n5278), 
	.A1(\fifo_from_fir/fifo_cell10/data_out/N35 ), 
	.A0(FE_OFN546_n4705));
   NOR2X1TS U5330 (.Y(n4526), 
	.B(FE_OFN223_n4525), 
	.A(FE_OFN840_n7619));
   AOI31X1TS U5331 (.Y(n4476), 
	.B0(\fifo_from_fft/hold[9] ), 
	.A2(n5318), 
	.A1(\fifo_from_fft/fifo_cell9/data_out/N35 ), 
	.A0(n4525));
   NOR2X1TS U5332 (.Y(n4712), 
	.B(FE_OFN560_n4711), 
	.A(FE_OFN837_n7619));
   AOI31X1TS U5333 (.Y(n4662), 
	.B0(\fifo_from_fir/hold[9] ), 
	.A2(n5279), 
	.A1(\fifo_from_fir/fifo_cell9/data_out/N35 ), 
	.A0(n4711));
   NOR2X1TS U5338 (.Y(n4532), 
	.B(FE_OFN233_n4531), 
	.A(FE_OFN840_n7619));
   NOR3X1TS U5339 (.Y(n4531), 
	.C(n4623), 
	.B(n4622), 
	.A(n8838));
   NOR3X1TS U5340 (.Y(n4717), 
	.C(n4809), 
	.B(n4808), 
	.A(n8871));
   NOR2X1TS U5341 (.Y(n4538), 
	.B(FE_OFN247_n4537), 
	.A(FE_OFN847_n7619));
   AOI31X1TS U5342 (.Y(n4472), 
	.B0(\fifo_from_fft/hold[7] ), 
	.A2(n5320), 
	.A1(\fifo_from_fft/fifo_cell7/data_out/N35 ), 
	.A0(FE_OFN247_n4537));
   AOI31X1TS U5343 (.Y(n4658), 
	.B0(\fifo_from_fir/hold[7] ), 
	.A2(n5281), 
	.A1(\fifo_from_fir/fifo_cell7/data_out/N35 ), 
	.A0(FE_OFN593_n4723));
   NOR2X1TS U5344 (.Y(n4724), 
	.B(FE_OFN595_n4723), 
	.A(FE_OFN837_n7619));
   NOR3X1TS U5346 (.Y(n4537), 
	.C(n4626), 
	.B(n4625), 
	.A(n8838));
   NOR3X1TS U5348 (.Y(n4723), 
	.C(n4812), 
	.B(n4811), 
	.A(n8871));
   AOI31X1TS U5349 (.Y(n4470), 
	.B0(\fifo_from_fft/hold[6] ), 
	.A2(n5321), 
	.A1(\fifo_from_fft/fifo_cell6/data_out/N35 ), 
	.A0(n4543));
   NOR2X1TS U5350 (.Y(n4544), 
	.B(FE_OFN267_n4543), 
	.A(FE_OFN835_n7619));
   AOI31X1TS U5351 (.Y(n4656), 
	.B0(\fifo_from_fir/hold[6] ), 
	.A2(n5282), 
	.A1(\fifo_from_fir/fifo_cell6/data_out/N35 ), 
	.A0(n4729));
   NOR3X1TS U5352 (.Y(n4543), 
	.C(n4629), 
	.B(n4628), 
	.A(n8838));
   NOR3X1TS U5353 (.Y(n4729), 
	.C(n4815), 
	.B(n4814), 
	.A(n8871));
   NOR2X1TS U5354 (.Y(n4550), 
	.B(FE_OFN290_n4549), 
	.A(FE_OFN844_n7619));
   AOI31X1TS U5355 (.Y(n4468), 
	.B0(\fifo_from_fft/hold[5] ), 
	.A2(n5322), 
	.A1(\fifo_from_fft/fifo_cell5/data_out/N35 ), 
	.A0(n4549));
   NOR2XLTS U5356 (.Y(n4736), 
	.B(FE_OFN621_n4735), 
	.A(FE_OFN845_n7619));
   AOI31X1TS U5357 (.Y(n4654), 
	.B0(\fifo_from_fir/hold[5] ), 
	.A2(n5283), 
	.A1(\fifo_from_fir/fifo_cell5/data_out/N35 ), 
	.A0(FE_OFN618_n4735));
   NOR3X1TS U5358 (.Y(n4549), 
	.C(n4632), 
	.B(n4631), 
	.A(n8837));
   AOI31X1TS U5359 (.Y(n4466), 
	.B0(\fifo_from_fft/hold[4] ), 
	.A2(n5323), 
	.A1(\fifo_from_fft/fifo_cell4/data_out/N35 ), 
	.A0(n4555));
   NOR2X1TS U5360 (.Y(n4556), 
	.B(FE_OFN302_n4555), 
	.A(FE_OFN835_n7619));
   AOI31X1TS U5361 (.Y(n4652), 
	.B0(\fifo_from_fir/hold[4] ), 
	.A2(n5284), 
	.A1(\fifo_from_fir/fifo_cell4/data_out/N35 ), 
	.A0(FE_OFN642_n4741));
   NOR2X1TS U5362 (.Y(n4742), 
	.B(FE_OFN646_n4741), 
	.A(FE_OFN845_n7619));
   NOR3X1TS U5363 (.Y(n4555), 
	.C(n4635), 
	.B(n4634), 
	.A(n8837));
   AOI31X1TS U5364 (.Y(n4464), 
	.B0(\fifo_from_fft/hold[3] ), 
	.A2(n5324), 
	.A1(\fifo_from_fft/fifo_cell3/data_out/N35 ), 
	.A0(FE_OFN313_n4561));
   AOI31X1TS U5365 (.Y(n4650), 
	.B0(\fifo_from_fir/hold[3] ), 
	.A2(n5285), 
	.A1(\fifo_from_fir/fifo_cell3/data_out/N35 ), 
	.A0(FE_OFN653_n4747));
   AOI31X1TS U5370 (.Y(n4648), 
	.B0(\fifo_from_fir/hold[2] ), 
	.A2(n5286), 
	.A1(\fifo_from_fir/fifo_cell2/data_out/N35 ), 
	.A0(n8137));
   NOR2X1TS U5371 (.Y(n3722), 
	.B(n3754), 
	.A(FE_OFN765_n3720));
   AOI21X1TS U5373 (.Y(n3531), 
	.B0(FE_OFN903_n3530), 
	.A1(n3564), 
	.A0(n3563));
   AOI21X1TS U5375 (.Y(n3575), 
	.B0(FE_OFN921_n3574), 
	.A1(n3608), 
	.A0(n3607));
   NOR2X1TS U5376 (.Y(n3721), 
	.B(n3755), 
	.A(n3720));
   AOI21X1TS U5377 (.Y(n3663), 
	.B0(FE_OFN881_n3662), 
	.A1(n3696), 
	.A0(n3695));
   AOI21X1TS U5378 (.Y(n3619), 
	.B0(FE_OFN970_n3618), 
	.A1(n3652), 
	.A0(n3651));
   OR3X1TS U5381 (.Y(n8056), 
	.C(n4641), 
	.B(n4640), 
	.A(n8837));
   AOI31X1TS U5383 (.Y(n4646), 
	.B0(\fifo_from_fir/hold[1] ), 
	.A2(n5287), 
	.A1(\fifo_from_fir/fifo_cell1/data_out/N35 ), 
	.A0(FE_OFN666_n4759));
   AOI31X1TS U5384 (.Y(n4460), 
	.B0(\fifo_from_fft/hold[1] ), 
	.A2(n5326), 
	.A1(\fifo_from_fft/fifo_cell1/data_out/N35 ), 
	.A0(n4573));
   NAND2X1TS U5385 (.Y(n3754), 
	.B(n3829), 
	.A(n7203));
   AOI21X1TS U5387 (.Y(n3487), 
	.B0(FE_OFN944_n3486), 
	.A1(n3520), 
	.A0(n3519));
   AND4X1TS U5388 (.Y(n8058), 
	.D(n3484), 
	.C(n9465), 
	.B(\router/fft_put_req_reg ), 
	.A(n3714));
   OA21XLTS U5392 (.Y(n4702), 
	.B0(n9486), 
	.A1(\fifo_from_fir/fifo_cell11/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell11/controller/f_i_get ));
   OA21XLTS U5393 (.Y(n4756), 
	.B0(n9484), 
	.A1(\fifo_from_fir/fifo_cell2/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell2/controller/f_i_get ));
   OA21XLTS U5394 (.Y(n4696), 
	.B0(n9487), 
	.A1(\fifo_from_fir/fifo_cell12/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell12/controller/f_i_get ));
   OA21XLTS U5395 (.Y(n4762), 
	.B0(n9484), 
	.A1(\fifo_from_fir/fifo_cell1/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell1/controller/f_i_get ));
   OA21XLTS U5396 (.Y(n4750), 
	.B0(n9484), 
	.A1(\fifo_from_fir/fifo_cell3/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell3/controller/f_i_get ));
   OA21XLTS U5397 (.Y(n4690), 
	.B0(n9487), 
	.A1(\fifo_from_fir/fifo_cell13/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell13/controller/f_i_get ));
   OA21XLTS U5398 (.Y(n4684), 
	.B0(n9487), 
	.A1(\fifo_from_fir/fifo_cell14/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell14/controller/f_i_get ));
   OA21XLTS U5399 (.Y(n4516), 
	.B0(n9482), 
	.A1(\fifo_from_fft/fifo_cell11/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell11/controller/f_i_get ));
   OA21XLTS U5400 (.Y(n4558), 
	.B0(n9480), 
	.A1(\fifo_from_fft/fifo_cell4/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell4/controller/f_i_get ));
   OA21XLTS U5401 (.Y(n4528), 
	.B0(n9482), 
	.A1(\fifo_from_fft/fifo_cell9/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell9/controller/f_i_get ));
   OA21XLTS U5402 (.Y(n4708), 
	.B0(n9486), 
	.A1(\fifo_from_fir/fifo_cell10/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell10/controller/f_i_get ));
   OA21XLTS U5403 (.Y(n4522), 
	.B0(n9482), 
	.A1(\fifo_from_fft/fifo_cell10/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell10/controller/f_i_get ));
   OA21XLTS U5404 (.Y(n4714), 
	.B0(n9486), 
	.A1(\fifo_from_fir/fifo_cell9/controller/f_i_put ), 
	.A0(\fifo_from_fir/fifo_cell9/controller/f_i_get ));
   INVX2TS U5405 (.Y(n9485), 
	.A(FE_OFN829_n7619));
   OA21XLTS U5406 (.Y(n4576), 
	.B0(n9497), 
	.A1(\fifo_from_fft/fifo_cell1/controller/f_i_put ), 
	.A0(\fifo_from_fft/fifo_cell1/controller/f_i_get ));
   AOI211X1TS U5407 (.Y(n3715), 
	.C0(n3713), 
	.B0(n9432), 
	.A1(n7953), 
	.A0(n9406));
   NAND3X1TS U5408 (.Y(n3713), 
	.C(n7211), 
	.B(n3850), 
	.A(n9407));
   NOR4XLTS U5410 (.Y(n3563), 
	.D(n3572), 
	.C(n3571), 
	.B(n3570), 
	.A(n3569));
   NOR4XLTS U5411 (.Y(n3519), 
	.D(n3528), 
	.C(n3527), 
	.B(n3526), 
	.A(n3525));
   NOR4XLTS U5412 (.Y(n3607), 
	.D(n3616), 
	.C(n3615), 
	.B(n3614), 
	.A(n3613));
   NOR4XLTS U5413 (.Y(n3695), 
	.D(n3704), 
	.C(n3703), 
	.B(n3702), 
	.A(n3701));
   NOR4XLTS U5414 (.Y(n3651), 
	.D(n3660), 
	.C(n3659), 
	.B(n3658), 
	.A(n3657));
   NOR4XLTS U5415 (.Y(n3608), 
	.D(n3612), 
	.C(n3611), 
	.B(n3610), 
	.A(n3609));
   NOR4XLTS U5416 (.Y(n3564), 
	.D(n3568), 
	.C(n3567), 
	.B(n3566), 
	.A(n3565));
   NOR4XLTS U5417 (.Y(n3652), 
	.D(n3656), 
	.C(n3655), 
	.B(n3654), 
	.A(n3653));
   NOR4XLTS U5418 (.Y(n3696), 
	.D(n3700), 
	.C(n3699), 
	.B(n3698), 
	.A(n3697));
   NOR4XLTS U5419 (.Y(n3520), 
	.D(n3524), 
	.C(n3523), 
	.B(n3522), 
	.A(n3521));
   NOR3X1TS U5420 (.Y(n6768), 
	.C(\fifo_to_fft/fifo_cell7/controller/write_enable ), 
	.B(n7301), 
	.A(\fifo_to_fft/fifo_cell7/controller/valid_read ));
   AOI31X1TS U5421 (.Y(n3865), 
	.B0(\fifo_to_fft/hold[7] ), 
	.A2(n6768), 
	.A1(\fifo_to_fft/fifo_cell7/data_out/N35 ), 
	.A0(n3927));
   NOR3X1TS U5422 (.Y(n6769), 
	.C(\fifo_to_fft/fifo_cell10/controller/write_enable ), 
	.B(n7276), 
	.A(\fifo_to_fft/fifo_cell10/controller/valid_read ));
   AOI31X1TS U5423 (.Y(n3871), 
	.B0(\fifo_to_fft/hold[10] ), 
	.A2(n6769), 
	.A1(\fifo_to_fft/fifo_cell10/data_out/N35 ), 
	.A0(n3912));
   CLKINVX1TS U5424 (.Y(n6770), 
	.A(n4067));
   AOI2BB2X1TS U5425 (.Y(n6771), 
	.B1(n6770), 
	.B0(n7366), 
	.A1N(n7365), 
	.A0N(n6770));
   AOI2BB2X1TS U5426 (.Y(n6772), 
	.B1(n7394), 
	.B0(n7404), 
	.A1N(n7395), 
	.A0N(n7405));
   XOR2X1TS U5427 (.Y(n6773), 
	.B(n4198), 
	.A(n6772));
   XOR2X1TS U5428 (.Y(n6774), 
	.B(n4127), 
	.A(n4122));
   XOR2X1TS U5429 (.Y(n6775), 
	.B(n6774), 
	.A(n6773));
   XOR2X1TS U5430 (.Y(n6776), 
	.B(n6775), 
	.A(n4087));
   CLKINVX1TS U5431 (.Y(n6777), 
	.A(n4107));
   AOI2BB2X1TS U5432 (.Y(n6778), 
	.B1(n6777), 
	.B0(n7425), 
	.A1N(n7424), 
	.A0N(n6777));
   XOR2X1TS U5433 (.Y(n6779), 
	.B(n6778), 
	.A(n4117));
   XOR2X1TS U5434 (.Y(n6780), 
	.B(n6779), 
	.A(n6776));
   XOR2X1TS U5435 (.Y(n6781), 
	.B(n6780), 
	.A(n6771));
   CLKINVX1TS U5436 (.Y(n6782), 
	.A(n4082));
   AOI2BB2X1TS U5437 (.Y(n6783), 
	.B1(n6782), 
	.B0(n7375), 
	.A1N(n7374), 
	.A0N(n6782));
   XOR2X1TS U5438 (.Y(n6784), 
	.B(n4102), 
	.A(n6783));
   XOR2X1TS U5439 (.Y(n6785), 
	.B(n6784), 
	.A(n6781));
   XOR2X1TS U5440 (.Y(n3804), 
	.B(n4062), 
	.A(n6785));
   NOR4XLTS U5441 (.Y(n6786), 
	.D(\fifo_to_fft/fifo_cell15/controller/write_enable ), 
	.C(n7242), 
	.B(n7236), 
	.A(n3881));
   CLKINVX1TS U5442 (.Y(n6787), 
	.A(\fifo_to_fft/fifo_cell15/controller/valid_read ));
   AO21X1TS U5443 (.Y(n3880), 
	.B0(\fifo_to_fft/hold[15] ), 
	.A1(n6787), 
	.A0(n6786));
   AOI222XLTS U5444 (.Y(n3733), 
	.C1(fir_data_in[20]), 
	.C0(FE_OFN752_n3722), 
	.B1(fft_data_in[20]), 
	.B0(FE_OFN762_n3721), 
	.A1(\router/data_cntl/data_in[20] ), 
	.A0(FE_OFN773_n3720));
   AOI222XLTS U5445 (.Y(n3726), 
	.C1(fir_data_in[27]), 
	.C0(FE_OFN747_n3722), 
	.B1(FE_MDBN10_), 
	.B0(FE_OFN757_n3721), 
	.A1(\router/data_cntl/data_in[27] ), 
	.A0(FE_OFN768_n3720));
   NOR3X1TS U5446 (.Y(n6788), 
	.C(\fifo_from_fft/fifo_cell2/controller/write_enable ), 
	.B(n7519), 
	.A(\fifo_from_fft/fifo_cell2/controller/valid_read ));
   AOI31X1TS U5447 (.Y(n4462), 
	.B0(\fifo_from_fft/hold[2] ), 
	.A2(n6788), 
	.A1(\fifo_from_fft/fifo_cell2/data_out/N35 ), 
	.A0(n8472));
   NOR3X1TS U5448 (.Y(n6789), 
	.C(\fifo_to_fir/fifo_cell2/controller/write_enable ), 
	.B(n7440), 
	.A(\fifo_to_fir/fifo_cell2/controller/valid_read ));
   AOI31X1TS U5449 (.Y(n4030), 
	.B0(\fifo_to_fir/hold[2] ), 
	.A2(n6789), 
	.A1(\fifo_to_fir/fifo_cell2/data_out/N35 ), 
	.A0(n4127));
   NOR3X1TS U5450 (.Y(n6790), 
	.C(\fifo_to_fir/fifo_cell6/controller/write_enable ), 
	.B(n7415), 
	.A(\fifo_to_fir/fifo_cell6/controller/valid_read ));
   AOI31X1TS U5451 (.Y(n4038), 
	.B0(\fifo_to_fir/hold[6] ), 
	.A2(n6790), 
	.A1(\fifo_to_fir/fifo_cell6/data_out/N35 ), 
	.A0(n4107));
   NOR3X1TS U5452 (.Y(n6791), 
	.C(\fifo_to_fir/fifo_cell11/controller/write_enable ), 
	.B(n7380), 
	.A(\fifo_to_fir/fifo_cell11/controller/valid_read ));
   AOI31X1TS U5453 (.Y(n4048), 
	.B0(\fifo_to_fir/hold[11] ), 
	.A2(n6791), 
	.A1(\fifo_to_fir/fifo_cell11/data_out/N35 ), 
	.A0(n4082));
   NAND2X1TS U5454 (.Y(n6792), 
	.B(n9515), 
	.A(n5288));
   OAI31X1TS U5455 (.Y(n3767), 
	.B0(\fifo_from_fir/fifo_cell0/reg_ptok/N29 ), 
	.A2(n6792), 
	.A1(\fifo_from_fir/fifo_cell0/reg_ptok/out_valid_put ), 
	.A0(\fifo_from_fir/fifo_cell0/reg_ptok/out_valid_get ));
   CLKINVX1TS U5456 (.Y(n6793), 
	.A(n3907));
   AOI2BB2X1TS U5457 (.Y(n6794), 
	.B1(n6793), 
	.B0(n7266), 
	.A1N(n7265), 
	.A0N(n6793));
   CLKINVX1TS U5458 (.Y(n6795), 
	.A(n3932));
   AOI2BB2X1TS U5459 (.Y(n6796), 
	.B1(n6795), 
	.B0(n7316), 
	.A1N(n7315), 
	.A0N(n6795));
   AOI2BB2X1TS U5460 (.Y(n6797), 
	.B1(n7285), 
	.B0(FE_OFN678_n7295), 
	.A1N(n7286), 
	.A0N(FE_OFN678_n7295));
   XOR2X1TS U5461 (.Y(n6798), 
	.B(n4023), 
	.A(n6797));
   XOR2X1TS U5462 (.Y(n6799), 
	.B(n3952), 
	.A(n3947));
   XOR2X1TS U5463 (.Y(n6800), 
	.B(n6799), 
	.A(n6798));
   XOR2X1TS U5464 (.Y(n6801), 
	.B(n6800), 
	.A(n3912));
   XOR2X1TS U5465 (.Y(n6802), 
	.B(n6796), 
	.A(n3942));
   XOR2X1TS U5466 (.Y(n6803), 
	.B(n6802), 
	.A(n6801));
   CLKINVX1TS U5467 (.Y(n6804), 
	.A(n3892));
   AOI2BB2X1TS U5468 (.Y(n6805), 
	.B1(n6804), 
	.B0(n7256), 
	.A1N(n7255), 
	.A0N(n6804));
   XOR2X1TS U5469 (.Y(n6806), 
	.B(n6803), 
	.A(n6805));
   XOR2X1TS U5470 (.Y(n6807), 
	.B(n3927), 
	.A(n6794));
   XOR2X1TS U5471 (.Y(n6808), 
	.B(n6807), 
	.A(n6806));
   XOR2X1TS U5472 (.Y(n3815), 
	.B(n3887), 
	.A(n6808));
   NOR4XLTS U5473 (.Y(n6809), 
	.D(\fifo_to_fir/fifo_cell15/controller/write_enable ), 
	.C(n7351), 
	.B(n7345), 
	.A(n4056));
   CLKINVX1TS U5474 (.Y(n6810), 
	.A(\fifo_to_fir/fifo_cell15/controller/valid_read ));
   AO21X1TS U5475 (.Y(n4055), 
	.B0(\fifo_to_fir/hold[15] ), 
	.A1(n6810), 
	.A0(n6809));
   NOR4X1TS U5476 (.Y(n6811), 
	.D(n7241), 
	.C(n7246), 
	.B(n7251), 
	.A(n7260));
   NOR4X1TS U5477 (.Y(n6812), 
	.D(n7270), 
	.C(n7275), 
	.B(n7280), 
	.A(n7290));
   NOR4X1TS U5478 (.Y(n6813), 
	.D(n7300), 
	.C(n7305), 
	.B(n7310), 
	.A(n7320));
   NOR4X1TS U5479 (.Y(n6814), 
	.D(n7325), 
	.C(n7330), 
	.B(n7340), 
	.A(n7231));
   NAND4X2TS U5480 (.Y(n3484), 
	.D(n6814), 
	.C(n6813), 
	.B(n6812), 
	.A(n6811));
   NOR4X1TS U5481 (.Y(n6815), 
	.D(n7528), 
	.C(n7533), 
	.B(n7538), 
	.A(n7543));
   NOR4X1TS U5482 (.Y(n6816), 
	.D(n7548), 
	.C(n7553), 
	.B(n7558), 
	.A(n7563));
   NOR4X1TS U5483 (.Y(n6817), 
	.D(n7568), 
	.C(n7573), 
	.B(n7578), 
	.A(n7583));
   NOR4XLTS U5484 (.Y(n6818), 
	.D(n7588), 
	.C(n7593), 
	.B(n7598), 
	.A(n7216));
   NAND4X2TS U5485 (.Y(n3465), 
	.D(n6818), 
	.C(n6817), 
	.B(n6816), 
	.A(n6815));
   NOR2X1TS U5486 (.Y(n6819), 
	.B(n3784), 
	.A(n3783));
   OAI2BB2XLTS U5487 (.Y(n6820), 
	.B1(FE_OFN783_n7619), 
	.B0(FE_OFN698_n8052), 
	.A1N(n6819), 
	.A0N(n3787));
   OAI211X1TS U5488 (.Y(n5418), 
	.C0(n6820), 
	.B0(n9464), 
	.A1(n3780), 
	.A0(FE_OFN698_n8052));
   AOI222XLTS U5489 (.Y(n3734), 
	.C1(fir_data_in[19]), 
	.C0(FE_OFN750_n3722), 
	.B1(fft_data_in[19]), 
	.B0(FE_OFN760_n3721), 
	.A1(\router/data_cntl/data_in[19] ), 
	.A0(FE_OFN771_n3720));
   AOI222XLTS U5490 (.Y(n3725), 
	.C1(FE_MDBN0_), 
	.C0(FE_OFN746_n3722), 
	.B1(FE_MDBN11_), 
	.B0(FE_OFN755_n3721), 
	.A1(\router/data_cntl/data_in[28] ), 
	.A0(FE_OFN767_n3720));
   NOR2BX1TS U5491 (.Y(\add_x_22_1/carry[31] ), 
	.B(n7367), 
	.AN(\add_x_22_1/carry[30] ));
   XNOR2X1TS U5492 (.Y(\router/addr_calc/fft_write_calc/counter/N76 ), 
	.B(\add_x_22_1/carry[30] ), 
	.A(n7367));
   NOR2BX1TS U5493 (.Y(\add_x_22_0/carry[30] ), 
	.B(n7491), 
	.AN(\add_x_22_0/carry[29] ));
   XNOR2X1TS U5494 (.Y(\router/addr_calc/fft_read_calc/counter/N75 ), 
	.B(\add_x_22_0/carry[29] ), 
	.A(n7491));
   NOR2BX1TS U5495 (.Y(\add_x_22_3/carry[30] ), 
	.B(n7123), 
	.AN(\add_x_22_3/carry[29] ));
   XNOR2X1TS U5496 (.Y(\router/addr_calc/fir_write_calc/counter/N75 ), 
	.B(\add_x_22_3/carry[29] ), 
	.A(n7123));
   NAND3X1TS U5497 (.Y(n6821), 
	.C(n7309), 
	.B(FE_OFN1271_router_addr_calc_fir_read_calc_count_15_), 
	.A(n7304));
   NAND4X1TS U5498 (.Y(n6822), 
	.D(n7359), 
	.C(n7354), 
	.B(n7364), 
	.A(\router/addr_calc/fir_read_calc/count[0] ));
   AND4X1TS U5499 (.Y(n6823), 
	.D(n7349), 
	.C(n7344), 
	.B(n7339), 
	.A(FE_OFN1276_router_addr_calc_fir_read_calc_count_5_));
   NAND4X1TS U5500 (.Y(n6824), 
	.D(n6823), 
	.C(n7329), 
	.B(n7334), 
	.A(\router/addr_calc/fir_read_calc/count[9] ));
   NAND3X1TS U5501 (.Y(n6825), 
	.C(n7314), 
	.B(n7319), 
	.A(n7324));
   NAND3X1TS U5502 (.Y(n6826), 
	.C(FE_OFN1260_router_addr_calc_fir_read_calc_count_19_), 
	.B(n7299), 
	.A(n7294));
   NOR4XLTS U5503 (.Y(n6827), 
	.D(n6826), 
	.C(n6825), 
	.B(n6824), 
	.A(n6822));
   NAND4X1TS U5504 (.Y(n6828), 
	.D(n6827), 
	.C(n7289), 
	.B(FE_OFN1250_n7278), 
	.A(FE_OFN1253_n7283));
   NAND3X1TS U5505 (.Y(n6829), 
	.C(FE_OFN1242_n7268), 
	.B(FE_OFN1243_n7273), 
	.A(FE_OFN1247_router_addr_calc_fir_read_calc_count_23_));
   NAND3X1TS U5506 (.Y(n6830), 
	.C(n7258), 
	.B(n7263), 
	.A(\router/addr_calc/fir_read_calc/count[27] ));
   NOR4XLTS U5507 (.Y(n6831), 
	.D(n6830), 
	.C(n6829), 
	.B(n6828), 
	.A(n6821));
   NAND4X1TS U5508 (.Y(\router/addr_calc/fir_read_calc/counter/N40 ), 
	.D(FE_OFN1230_router_addr_calc_fir_read_calc_count_30_), 
	.C(n7249), 
	.B(FE_OFN1235_n7254), 
	.A(n6831));
   NOR3X1TS U5509 (.Y(n6832), 
	.C(\fifo_to_fft/fifo_cell3/controller/write_enable ), 
	.B(n7326), 
	.A(\fifo_to_fft/fifo_cell3/controller/valid_read ));
   AOI31X1TS U5510 (.Y(n3857), 
	.B0(\fifo_to_fft/hold[3] ), 
	.A2(n6832), 
	.A1(\fifo_to_fft/fifo_cell3/data_out/N35 ), 
	.A0(n3947));
   NOR3X1TS U5511 (.Y(n6833), 
	.C(\fifo_to_fft/fifo_cell6/controller/write_enable ), 
	.B(n7306), 
	.A(\fifo_to_fft/fifo_cell6/controller/valid_read ));
   AOI31X1TS U5512 (.Y(n3863), 
	.B0(\fifo_to_fft/hold[6] ), 
	.A2(n6833), 
	.A1(\fifo_to_fft/fifo_cell6/data_out/N35 ), 
	.A0(n3932));
   NOR3X1TS U5513 (.Y(n6834), 
	.C(\fifo_to_fft/fifo_cell9/controller/write_enable ), 
	.B(n7281), 
	.A(\fifo_to_fft/fifo_cell9/controller/valid_read ));
   AOI31X1TS U5514 (.Y(n3869), 
	.B0(\fifo_to_fft/hold[9] ), 
	.A2(n6834), 
	.A1(\fifo_to_fft/fifo_cell9/data_out/N35 ), 
	.A0(n7285));
   XOR2X1TS U5515 (.Y(n6835), 
	.B(FE_OFN555_n4705), 
	.A(FE_OFN474_n4675));
   AOI2BB2X1TS U5516 (.Y(n6836), 
	.B1(FE_OFN511_n4693), 
	.B0(FE_OFN543_n4699), 
	.A1N(FE_OFN511_n4693), 
	.A0N(FE_OFN543_n4699));
   XOR2XLTS U5517 (.Y(n6837), 
	.B(n4781), 
	.A(FE_OFN641_n4741));
   XOR2X1TS U5518 (.Y(n6838), 
	.B(n8053), 
	.A(FE_OFN652_n4747));
   XOR2X1TS U5519 (.Y(n6839), 
	.B(n6838), 
	.A(n6837));
   XOR2XLTS U5520 (.Y(n6840), 
	.B(n6839), 
	.A(FE_OFN568_n4711));
   AOI2BB2X1TS U5521 (.Y(n6841), 
	.B1(FE_OFN580_n4717), 
	.B0(FE_OFN602_n4723), 
	.A1N(FE_OFN580_n4717), 
	.A0N(FE_OFN602_n4723));
   AOI2BB2X1TS U5522 (.Y(n6842), 
	.B1(FE_OFN612_n4729), 
	.B0(FE_OFN626_n4735), 
	.A1N(FE_OFN612_n4729), 
	.A0N(FE_OFN626_n4735));
   XOR2X1TS U5523 (.Y(n6843), 
	.B(n6842), 
	.A(n6841));
   XOR2X1TS U5524 (.Y(n6844), 
	.B(n6843), 
	.A(n6840));
   XOR2X1TS U5525 (.Y(n6845), 
	.B(n6844), 
	.A(n6836));
   XOR2X1TS U5526 (.Y(n6846), 
	.B(n6845), 
	.A(n6835));
   CLKINVX1TS U5527 (.Y(n6847), 
	.A(FE_OFN508_n8055));
   AOI2BB2X1TS U5528 (.Y(n6848), 
	.B1(n6847), 
	.B0(n4681), 
	.A1N(FE_OFN497_n4681), 
	.A0N(n6847));
   XOR2X1TS U5529 (.Y(n3764), 
	.B(n6848), 
	.A(n6846));
   NOR3X1TS U5530 (.Y(n6849), 
	.C(\fifo_to_fft/fifo_cell12/controller/write_enable ), 
	.B(n7261), 
	.A(\fifo_to_fft/fifo_cell12/controller/valid_read ));
   AOI31X1TS U5531 (.Y(n3875), 
	.B0(\fifo_to_fft/hold[12] ), 
	.A2(n6849), 
	.A1(\fifo_to_fft/fifo_cell12/data_out/N35 ), 
	.A0(n7265));
   NAND2X1TS U5532 (.Y(n6850), 
	.B(n9515), 
	.A(n5327));
   OAI31X1TS U5533 (.Y(n3787), 
	.B0(\fifo_from_fft/fifo_cell0/reg_ptok/N29 ), 
	.A2(n6850), 
	.A1(\fifo_from_fft/fifo_cell0/reg_ptok/out_valid_put ), 
	.A0(\fifo_from_fft/fifo_cell0/reg_ptok/out_valid_get ));
   NOR3X1TS U5534 (.Y(n6851), 
	.C(\fifo_to_fft/fifo_cell14/controller/write_enable ), 
	.B(n7247), 
	.A(\fifo_to_fft/fifo_cell14/controller/valid_read ));
   AOI31X1TS U5535 (.Y(n3879), 
	.B0(\fifo_to_fft/hold[14] ), 
	.A2(n6851), 
	.A1(n3892), 
	.A0(\fifo_to_fft/fifo_cell14/data_out/N35 ));
   NOR4X1TS U5536 (.Y(n6852), 
	.D(n7162), 
	.C(FE_OFN1244_router_addr_calc_iir_write_calc_count_23_), 
	.B(n7168), 
	.A(n7174));
   NAND2X1TS U5537 (.Y(n6853), 
	.B(n7113), 
	.A(n7952));
   NOR4XLTS U5538 (.Y(n6854), 
	.D(n7139), 
	.C(n7127), 
	.B(n7133), 
	.A(FE_OFN1441_router_addr_calc_iir_write_calc_count_16_));
   NOR4XLTS U5539 (.Y(n6855), 
	.D(n7151), 
	.C(n7157), 
	.B(n7145), 
	.A(FE_OFN1440_router_addr_calc_iir_write_calc_count_19_));
   NOR4XLTS U5540 (.Y(n6856), 
	.D(n7099), 
	.C(n7090), 
	.B(n7093), 
	.A(FE_OFN1280_router_addr_calc_iir_write_calc_count_9_));
   NOR4XLTS U5541 (.Y(n6857), 
	.D(n7116), 
	.C(n7122), 
	.B(n7105), 
	.A(n7110));
   NAND4X1TS U5542 (.Y(n6858), 
	.D(n6857), 
	.C(n6856), 
	.B(n6855), 
	.A(n6854));
   NOR4XLTS U5543 (.Y(n6859), 
	.D(n6858), 
	.C(n6853), 
	.B(n7180), 
	.A(FE_OFN1439_router_addr_calc_iir_write_calc_count_27_));
   OR4X1TS U5544 (.Y(n6860), 
	.D(n7106), 
	.C(n7186), 
	.B(n7198), 
	.A(FE_OFN1442_router_addr_calc_iir_write_calc_count_0_));
   NOR4XLTS U5545 (.Y(n6861), 
	.D(n6860), 
	.C(n7192), 
	.B(n7096), 
	.A(FE_OFN1281_router_addr_calc_iir_write_calc_count_5_));
   NAND4X1TS U5546 (.Y(\router/addr_calc/iir_write_calc/counter/N40 ), 
	.D(n6861), 
	.C(n7102), 
	.B(n6859), 
	.A(n6852));
   NOR4XLTS U5547 (.Y(n6862), 
	.D(n7454), 
	.C(n7459), 
	.B(n7464), 
	.A(n7469));
   NOR4X1TS U5548 (.Y(n6863), 
	.D(n7474), 
	.C(n7479), 
	.B(n7484), 
	.A(n7489));
   NOR4X1TS U5549 (.Y(n6864), 
	.D(n7493), 
	.C(n7498), 
	.B(n7503), 
	.A(n7508));
   NOR4X1TS U5550 (.Y(n6865), 
	.D(n7513), 
	.C(n7518), 
	.B(n7523), 
	.A(n7221));
   NAND4X2TS U5551 (.Y(n3477), 
	.D(n6865), 
	.C(n6864), 
	.B(n6863), 
	.A(n6862));
   NOR2BX1TS U5552 (.Y(n4136), 
	.B(n4181), 
	.AN(FE_OFN733_n8057));
   NOR4X1TS U5553 (.Y(n6866), 
	.D(n7350), 
	.C(n7355), 
	.B(n7360), 
	.A(n7369));
   NOR4XLTS U5554 (.Y(n6867), 
	.D(n7379), 
	.C(n7384), 
	.B(n7389), 
	.A(n7399));
   NOR4XLTS U5555 (.Y(n6868), 
	.D(n7409), 
	.C(n7414), 
	.B(n7419), 
	.A(n7429));
   NOR4XLTS U5556 (.Y(n6869), 
	.D(n7434), 
	.C(n7439), 
	.B(n7449), 
	.A(n7226));
   AND4X2TS U5557 (.Y(n3474), 
	.D(n6869), 
	.C(n6868), 
	.B(n6867), 
	.A(n6866));
   NOR4XLTS U5558 (.Y(n6870), 
	.D(\router/addr_calc/iir_read_calc/count[24] ), 
	.C(\router/addr_calc/iir_read_calc/count[25] ), 
	.B(\router/addr_calc/iir_read_calc/count[23] ), 
	.A(\router/addr_calc/iir_read_calc/count[22] ));
   NOR4XLTS U5559 (.Y(n6871), 
	.D(\router/addr_calc/iir_read_calc/count[29] ), 
	.C(\router/addr_calc/iir_read_calc/count[28] ), 
	.B(\router/addr_calc/iir_read_calc/count[0] ), 
	.A(\router/addr_calc/iir_read_calc/count[31] ));
   NOR4XLTS U5560 (.Y(n6872), 
	.D(\router/addr_calc/iir_read_calc/count[10] ), 
	.C(\router/addr_calc/iir_read_calc/count[13] ), 
	.B(\router/addr_calc/iir_read_calc/count[11] ), 
	.A(\router/addr_calc/iir_read_calc/count[12] ));
   NOR4XLTS U5561 (.Y(n6873), 
	.D(\router/addr_calc/iir_read_calc/count[8] ), 
	.C(\router/addr_calc/iir_read_calc/count[9] ), 
	.B(\router/addr_calc/iir_read_calc/count[7] ), 
	.A(\router/addr_calc/iir_read_calc/count[6] ));
   NAND4X1TS U5562 (.Y(n6874), 
	.D(n6873), 
	.C(n6872), 
	.B(n6871), 
	.A(\router/addr_calc/iir_read_calc/count[2] ));
   NOR3X1TS U5563 (.Y(n6875), 
	.C(n6874), 
	.B(\router/addr_calc/iir_read_calc/count[5] ), 
	.A(\router/addr_calc/iir_read_calc/count[4] ));
   NOR4XLTS U5564 (.Y(n6876), 
	.D(\router/addr_calc/iir_read_calc/count[20] ), 
	.C(\router/addr_calc/iir_read_calc/count[21] ), 
	.B(\router/addr_calc/iir_read_calc/count[19] ), 
	.A(\router/addr_calc/iir_read_calc/count[18] ));
   NOR4XLTS U5565 (.Y(n6877), 
	.D(\router/addr_calc/iir_read_calc/count[16] ), 
	.C(\router/addr_calc/iir_read_calc/count[17] ), 
	.B(\router/addr_calc/iir_read_calc/count[15] ), 
	.A(\router/addr_calc/iir_read_calc/count[14] ));
   NAND4X1TS U5566 (.Y(n6878), 
	.D(n6877), 
	.C(n6876), 
	.B(n6875), 
	.A(\router/addr_calc/iir_read_calc/count[3] ));
   NOR3X1TS U5567 (.Y(n6879), 
	.C(n6878), 
	.B(\router/addr_calc/iir_read_calc/count[27] ), 
	.A(\router/addr_calc/iir_read_calc/count[26] ));
   NAND4X1TS U5568 (.Y(\router/addr_calc/iir_read_calc/counter/N40 ), 
	.D(n6879), 
	.C(n6870), 
	.B(n8011), 
	.A(\router/addr_calc/iir_read_calc/count[1] ));
   NOR2X1TS U5569 (.Y(n6880), 
	.B(n3815), 
	.A(n3814));
   OAI2BB2XLTS U5570 (.Y(n6881), 
	.B1(FE_OFN782_n7619), 
	.B0(n8058), 
	.A1N(n6880), 
	.A0N(n3818));
   OAI211X1TS U5571 (.Y(n5455), 
	.C0(n6881), 
	.B0(n9463), 
	.A1(n3811), 
	.A0(n8058));
   NAND4X1TS U5572 (.Y(n6882), 
	.D(n7573), 
	.C(n7568), 
	.B(n7583), 
	.A(n7578));
   NAND4X1TS U5573 (.Y(n6883), 
	.D(n7598), 
	.C(n7593), 
	.B(n7588), 
	.A(n7216));
   NAND4X1TS U5574 (.Y(n6884), 
	.D(n7543), 
	.C(n7528), 
	.B(n7538), 
	.A(n7533));
   NAND4X1TS U5575 (.Y(n6885), 
	.D(n7553), 
	.C(n7563), 
	.B(n7558), 
	.A(n7548));
   NOR4X1TS U5576 (.Y(\fifo_from_fir/empty_det/N4 ), 
	.D(n6885), 
	.C(n6884), 
	.B(n6883), 
	.A(n6882));
   OAI21X1TS U5577 (.Y(n6886), 
	.B0(n4830), 
	.A1(\router/fir_get_req_reg ), 
	.A0(\router/iir_get_req_reg ));
   OAI2BB1X1TS U5578 (.Y(n6887), 
	.B0(n6886), 
	.A1N(FE_OFN1282_router_fft_get_req_reg), 
	.A0N(n7610));
   NOR3BX1TS U5579 (.Y(n6888), 
	.C(FE_OFN1282_router_fft_get_req_reg), 
	.B(FE_OFN990_n9431), 
	.AN(\router/fir_get_req_reg ));
   OAI21X1TS U5580 (.Y(n6889), 
	.B0(n7611), 
	.A1(n4832), 
	.A0(n9390));
   AOI211X1TS U5581 (.Y(n6890), 
	.C0(n6889), 
	.B0(n6888), 
	.A1(FE_OFN1282_router_fft_get_req_reg), 
	.A0(n9432));
   NAND4X1TS U5582 (.Y(n6891), 
	.D(n3832), 
	.C(n4644), 
	.B(n3754), 
	.A(n6890));
   CLKMX2X2TS U5583 (.Y(n6763), 
	.S0(n6891), 
	.B(n6887), 
	.A(\router/ram_write_enable_reg ));
   AOI222XLTS U5584 (.Y(n3746), 
	.C1(fir_data_in[7]), 
	.C0(FE_OFN745_n3722), 
	.B1(FE_MDBN15_), 
	.B0(FE_OFN756_n3721), 
	.A1(\router/data_cntl/data_in[7] ), 
	.A0(FE_OFN766_n3720));
   AOI222XLTS U5585 (.Y(n3732), 
	.C1(fir_data_in[21]), 
	.C0(FE_OFN752_n3722), 
	.B1(fft_data_in[21]), 
	.B0(FE_OFN762_n3721), 
	.A1(\router/data_cntl/data_in[21] ), 
	.A0(FE_OFN773_n3720));
   AOI222XLTS U5586 (.Y(n3724), 
	.C1(FE_MDBN1_), 
	.C0(n3722), 
	.B1(FE_MDBN12_), 
	.B0(FE_OFN755_n3721), 
	.A1(\router/data_cntl/data_in[29] ), 
	.A0(FE_OFN765_n3720));
   NAND4X1TS U5587 (.Y(n6892), 
	.D(instruction[26]), 
	.C(instruction[0]), 
	.B(instruction[29]), 
	.A(instruction[27]));
   NOR4XLTS U5588 (.Y(n6893), 
	.D(instruction[14]), 
	.C(instruction[15]), 
	.B(instruction[16]), 
	.A(instruction[17]));
   NOR4XLTS U5589 (.Y(n6894), 
	.D(instruction[10]), 
	.C(instruction[11]), 
	.B(instruction[12]), 
	.A(instruction[13]));
   NOR4XLTS U5590 (.Y(n6895), 
	.D(instruction[22]), 
	.C(instruction[23]), 
	.B(instruction[24]), 
	.A(instruction[25]));
   NOR4XLTS U5591 (.Y(n6896), 
	.D(instruction[18]), 
	.C(instruction[19]), 
	.B(instruction[20]), 
	.A(instruction[21]));
   NAND4X1TS U5592 (.Y(n6897), 
	.D(n6896), 
	.C(n6895), 
	.B(n6894), 
	.A(n6893));
   NOR3X1TS U5593 (.Y(n6898), 
	.C(n6897), 
	.B(n6892), 
	.A(n3458));
   NOR4BX1TS U5594 (.Y(n6899), 
	.D(instruction[7]), 
	.C(instruction[9]), 
	.B(instruction[8]), 
	.AN(instruction[28]));
   NOR4XLTS U5595 (.Y(n6900), 
	.D(instruction[3]), 
	.C(instruction[4]), 
	.B(instruction[5]), 
	.A(instruction[6]));
   NAND4X1TS U5596 (.Y(n4840), 
	.D(n6900), 
	.C(n6899), 
	.B(n6898), 
	.A(\router/pla_top/instruction_valid ));
   NAND3X1TS U5597 (.Y(n6901), 
	.C(n7547), 
	.B(n7542), 
	.A(FE_OFN1263_router_addr_calc_fft_read_calc_count_16_));
   NAND4X1TS U5598 (.Y(n6902), 
	.D(n7597), 
	.C(n7592), 
	.B(n7602), 
	.A(FE_OFN1444_router_addr_calc_fft_read_calc_count_0_));
   AND4X1TS U5599 (.Y(n6903), 
	.D(n7587), 
	.C(n7582), 
	.B(n7577), 
	.A(FE_OFN1273_router_addr_calc_fft_read_calc_count_5_));
   NAND4X1TS U5600 (.Y(n6904), 
	.D(n6903), 
	.C(n7567), 
	.B(n7572), 
	.A(FE_OFN1267_router_addr_calc_fft_read_calc_count_9_));
   NAND3X1TS U5601 (.Y(n6905), 
	.C(n7552), 
	.B(n7557), 
	.A(n7562));
   NAND3X1TS U5602 (.Y(n6906), 
	.C(FE_OFN1258_router_addr_calc_fft_read_calc_count_19_), 
	.B(n7537), 
	.A(n7532));
   NOR4XLTS U5603 (.Y(n6907), 
	.D(n6906), 
	.C(n6905), 
	.B(n6904), 
	.A(n6902));
   NAND4X1TS U5604 (.Y(n6908), 
	.D(n6907), 
	.C(n7527), 
	.B(n7516), 
	.A(n7521));
   NAND3X1TS U5605 (.Y(n6909), 
	.C(n7506), 
	.B(n7511), 
	.A(FE_OFN1245_router_addr_calc_fft_read_calc_count_23_));
   NAND3X1TS U5606 (.Y(n6910), 
	.C(n7496), 
	.B(n7501), 
	.A(FE_OFN1237_router_addr_calc_fft_read_calc_count_27_));
   NOR4X1TS U5607 (.Y(n6911), 
	.D(n6910), 
	.C(n6909), 
	.B(n6908), 
	.A(n6901));
   NAND4X1TS U5608 (.Y(\router/addr_calc/fft_read_calc/counter/N40 ), 
	.D(FE_OFN1229_router_addr_calc_fft_read_calc_count_30_), 
	.C(n7487), 
	.B(FE_OFN1234_n7492), 
	.A(n6911));
   NAND3X1TS U5609 (.Y(n6912), 
	.C(n7423), 
	.B(FE_OFN1270_router_addr_calc_fft_write_calc_count_15_), 
	.A(n7418));
   NAND4X1TS U5610 (.Y(n6913), 
	.D(n7478), 
	.C(n7473), 
	.B(n7483), 
	.A(\router/addr_calc/fft_write_calc/count[0] ));
   AND4X1TS U5611 (.Y(n6914), 
	.D(n7468), 
	.C(n7458), 
	.B(n7453), 
	.A(n7463));
   NAND4X1TS U5612 (.Y(n6915), 
	.D(n6914), 
	.C(n7443), 
	.B(n7448), 
	.A(\router/addr_calc/fft_write_calc/count[9] ));
   NAND3X1TS U5613 (.Y(n6916), 
	.C(n7428), 
	.B(n7433), 
	.A(n7438));
   NAND3X1TS U5614 (.Y(n6917), 
	.C(FE_OFN1259_router_addr_calc_fft_write_calc_count_19_), 
	.B(n7413), 
	.A(n7408));
   NOR4XLTS U5615 (.Y(n6918), 
	.D(n6917), 
	.C(n6916), 
	.B(n6915), 
	.A(n6913));
   NAND4X1TS U5616 (.Y(n6919), 
	.D(n6918), 
	.C(n7403), 
	.B(FE_OFN1249_n7392), 
	.A(FE_OFN1252_n7397));
   NAND3X1TS U5617 (.Y(n6920), 
	.C(n7382), 
	.B(n7387), 
	.A(FE_OFN1246_router_addr_calc_fft_write_calc_count_23_));
   NAND3X1TS U5618 (.Y(n6921), 
	.C(n7372), 
	.B(n7377), 
	.A(FE_OFN1238_router_addr_calc_fft_write_calc_count_27_));
   NOR4XLTS U5619 (.Y(n6922), 
	.D(n6921), 
	.C(n6920), 
	.B(n6919), 
	.A(n6912));
   NAND4X1TS U5620 (.Y(\router/addr_calc/fft_write_calc/counter/N40 ), 
	.D(FE_OFN1232_n7368), 
	.C(FE_OFN1228_router_addr_calc_fft_write_calc_count_31_), 
	.B(FE_OFN1233_router_addr_calc_fft_write_calc_count_29_), 
	.A(n6922));
   NAND3X1TS U5621 (.Y(n6923), 
	.C(n7190), 
	.B(n7184), 
	.A(FE_OFN1264_router_addr_calc_fir_write_calc_count_16_));
   NAND4X1TS U5622 (.Y(n6924), 
	.D(n7240), 
	.C(n7235), 
	.B(n7245), 
	.A(FE_OFN1445_router_addr_calc_fir_write_calc_count_0_));
   AND4X1TS U5623 (.Y(n6925), 
	.D(n7230), 
	.C(n7225), 
	.B(n7220), 
	.A(FE_OFN1272_router_addr_calc_fir_write_calc_count_5_));
   NAND4X1TS U5624 (.Y(n6926), 
	.D(n6925), 
	.C(n7210), 
	.B(n7215), 
	.A(\router/addr_calc/fir_write_calc/count[9] ));
   NAND3X1TS U5625 (.Y(n6927), 
	.C(n7196), 
	.B(n7202), 
	.A(n7206));
   NAND3X1TS U5626 (.Y(n6928), 
	.C(FE_OFN1261_router_addr_calc_fir_write_calc_count_19_), 
	.B(n7178), 
	.A(n7172));
   NOR4XLTS U5627 (.Y(n6929), 
	.D(n6928), 
	.C(n6927), 
	.B(n6926), 
	.A(n6924));
   NAND4X1TS U5628 (.Y(n6930), 
	.D(n6929), 
	.C(n7166), 
	.B(FE_OFN1251_n7153), 
	.A(FE_OFN1254_n7159));
   NAND3X1TS U5629 (.Y(n6931), 
	.C(n7141), 
	.B(n7147), 
	.A(\router/addr_calc/fir_write_calc/count[23] ));
   NAND3X1TS U5630 (.Y(n6932), 
	.C(n7129), 
	.B(n7135), 
	.A(FE_OFN1240_router_addr_calc_fir_write_calc_count_27_));
   NOR4XLTS U5631 (.Y(n6933), 
	.D(n6932), 
	.C(n6931), 
	.B(n6930), 
	.A(n6923));
   NAND4X1TS U5632 (.Y(\router/addr_calc/fir_write_calc/counter/N40 ), 
	.D(FE_OFN1231_router_addr_calc_fir_write_calc_count_30_), 
	.C(n7118), 
	.B(n7124), 
	.A(n6933));
   NOR3X1TS U5633 (.Y(n6934), 
	.C(\fifo_from_fir/fifo_cell8/controller/write_enable ), 
	.B(n7564), 
	.A(\fifo_from_fir/fifo_cell8/controller/valid_read ));
   AOI31X1TS U5634 (.Y(n4660), 
	.B0(\fifo_from_fir/hold[8] ), 
	.A2(n6934), 
	.A1(\fifo_from_fir/fifo_cell8/data_out/N35 ), 
	.A0(n4717));
   NOR3X1TS U5635 (.Y(n6935), 
	.C(\fifo_from_fir/fifo_cell15/controller/write_enable ), 
	.B(n7529), 
	.A(\fifo_from_fir/fifo_cell15/controller/valid_read ));
   AOI31X1TS U5636 (.Y(n4674), 
	.B0(\fifo_from_fir/hold[15] ), 
	.A2(n6935), 
	.A1(n4675), 
	.A0(\fifo_from_fir/fifo_cell15/data_out/N35 ));
   NOR2BX1TS U5637 (.Y(n3961), 
	.B(n4006), 
	.AN(n8058));
   AOI2BB2X1TS U5638 (.Y(n6936), 
	.B1(n4507), 
	.B0(n4513), 
	.A1N(n4507), 
	.A0N(n4513));
   AOI2BB2X1TS U5639 (.Y(n6937), 
	.B1(FE_OFN232_n4531), 
	.B0(FE_OFN250_n4537), 
	.A1N(FE_OFN232_n4531), 
	.A0N(FE_OFN250_n4537));
   AOI2BB2X1TS U5640 (.Y(n6938), 
	.B1(FE_OFN274_n4543), 
	.B0(FE_OFN289_n4549), 
	.A1N(FE_OFN274_n4543), 
	.A0N(FE_OFN289_n4549));
   XOR2X1TS U5641 (.Y(n6939), 
	.B(n4595), 
	.A(FE_OFN301_n4555));
   XOR2XLTS U5642 (.Y(n6940), 
	.B(n8056), 
	.A(FE_OFN320_n4561));
   XOR2X1TS U5643 (.Y(n6941), 
	.B(n6940), 
	.A(n6939));
   XOR2XLTS U5644 (.Y(n6942), 
	.B(n6941), 
	.A(n4525));
   XOR2X1TS U5645 (.Y(n6943), 
	.B(n6938), 
	.A(n6937));
   XOR2X1TS U5646 (.Y(n6944), 
	.B(n6943), 
	.A(n6942));
   XOR2X1TS U5647 (.Y(n6945), 
	.B(FE_OFN209_n4519), 
	.A(FE_OFN139_n4489));
   XOR2X1TS U5648 (.Y(n6946), 
	.B(n6944), 
	.A(n6936));
   XOR2X1TS U5649 (.Y(n6947), 
	.B(n6946), 
	.A(n6945));
   CLKINVX1TS U5650 (.Y(n6948), 
	.A(n8054));
   AOI2BB2X1TS U5651 (.Y(n6949), 
	.B1(n6948), 
	.B0(FE_OFN161_n4495), 
	.A1N(FE_OFN161_n4495), 
	.A0N(n6948));
   XOR2X1TS U5652 (.Y(n3784), 
	.B(n6949), 
	.A(n6947));
   NOR2X1TS U5653 (.Y(n6950), 
	.B(n3804), 
	.A(n3803));
   OAI2BB2XLTS U5654 (.Y(n6951), 
	.B1(FE_OFN787_n7619), 
	.B0(FE_OFN733_n8057), 
	.A1N(n6950), 
	.A0N(n3807));
   OAI211X1TS U5655 (.Y(n5453), 
	.C0(n6951), 
	.B0(n9463), 
	.A1(n3800), 
	.A0(FE_OFN732_n8057));
   NAND4X1TS U5656 (.Y(n6952), 
	.D(n7498), 
	.C(n7493), 
	.B(n7508), 
	.A(n7503));
   NAND4X1TS U5657 (.Y(n6953), 
	.D(n7523), 
	.C(n7518), 
	.B(n7513), 
	.A(n7221));
   NAND4X1TS U5658 (.Y(n6954), 
	.D(n7469), 
	.C(n7454), 
	.B(n7464), 
	.A(n7459));
   NAND4X1TS U5659 (.Y(n6955), 
	.D(n7479), 
	.C(n7489), 
	.B(n7484), 
	.A(n7474));
   NOR4XLTS U5660 (.Y(\fifo_from_fft/empty_det/N4 ), 
	.D(n6955), 
	.C(n6954), 
	.B(n6953), 
	.A(n6952));
   NAND4X1TS U5661 (.Y(n6956), 
	.D(n7414), 
	.C(n7409), 
	.B(n7429), 
	.A(n7419));
   NAND4X1TS U5662 (.Y(n6957), 
	.D(n7449), 
	.C(n7439), 
	.B(n7434), 
	.A(n7226));
   NAND4X1TS U5663 (.Y(n6958), 
	.D(n7369), 
	.C(n7350), 
	.B(n7360), 
	.A(n7355));
   NAND4X1TS U5664 (.Y(n6959), 
	.D(n7384), 
	.C(n7399), 
	.B(n7389), 
	.A(n7379));
   NOR4X1TS U5665 (.Y(\fifo_to_fir/empty_det/N4 ), 
	.D(n6959), 
	.C(n6958), 
	.B(n6957), 
	.A(n6956));
   NAND4X1TS U5666 (.Y(n6960), 
	.D(n7305), 
	.C(n7300), 
	.B(n7320), 
	.A(n7310));
   NAND4X1TS U5667 (.Y(n6961), 
	.D(n7340), 
	.C(n7330), 
	.B(n7325), 
	.A(n7231));
   NAND4X1TS U5668 (.Y(n6962), 
	.D(n7260), 
	.C(n7241), 
	.B(n7251), 
	.A(n7246));
   NAND4X1TS U5669 (.Y(n6963), 
	.D(n7275), 
	.C(n7290), 
	.B(n7280), 
	.A(n7270));
   NOR4X1TS U5670 (.Y(\fifo_to_fft/empty_det/N4 ), 
	.D(n6963), 
	.C(n6962), 
	.B(n6961), 
	.A(n6960));
   CLKINVX1TS U5671 (.Y(n6964), 
	.A(n4132));
   OAI211X1TS U5672 (.Y(n6965), 
	.C0(n9473), 
	.B0(\fifo_to_fir/hang[0] ), 
	.A1(n4026), 
	.A0(n8791));
   OAI31X1TS U5673 (.Y(n5569), 
	.B0(n6965), 
	.A2(n6964), 
	.A1(\fifo_to_fir/hang[0] ), 
	.A0(n4026));
   CLKINVX1TS U5674 (.Y(n6966), 
	.A(n3957));
   OAI211X1TS U5675 (.Y(n6967), 
	.C0(n9477), 
	.B0(\fifo_to_fft/hang[0] ), 
	.A1(n3851), 
	.A0(n8812));
   OAI31X1TS U5676 (.Y(n5517), 
	.B0(n6967), 
	.A2(n6966), 
	.A1(\fifo_to_fft/hang[0] ), 
	.A0(n3851));
   AOI222XLTS U5677 (.Y(n3753), 
	.C1(fir_data_in[0]), 
	.C0(FE_OFN746_n3722), 
	.B1(FE_MDBN3_), 
	.B0(FE_OFN756_n3721), 
	.A1(\router/data_cntl/data_in[0] ), 
	.A0(FE_OFN767_n3720));
   AOI222XLTS U5678 (.Y(n3731), 
	.C1(fir_data_in[22]), 
	.C0(FE_OFN752_n3722), 
	.B1(fft_data_in[22]), 
	.B0(FE_OFN762_n3721), 
	.A1(\router/data_cntl/data_in[22] ), 
	.A0(FE_OFN773_n3720));
   AOI222XLTS U5679 (.Y(n3723), 
	.C1(fir_data_in[30]), 
	.C0(FE_OFN745_n3722), 
	.B1(FE_MDBN13_), 
	.B0(FE_OFN756_n3721), 
	.A1(\router/data_cntl/data_in[30] ), 
	.A0(FE_OFN766_n3720));
   AOI22X1TS U5680 (.Y(n6968), 
	.B1(\fifo_from_fft/fifo_cell14/data_out/N35 ), 
	.B0(\fifo_from_fft/fifo_cell7/data_out/N35 ), 
	.A1(n4542), 
	.A0(n4500));
   AOI22X1TS U5681 (.Y(n6969), 
	.B1(\fifo_from_fft/fifo_cell12/data_out/N35 ), 
	.B0(\fifo_from_fft/fifo_cell11/data_out/N35 ), 
	.A1(n4512), 
	.A0(n4518));
   AOI22X1TS U5682 (.Y(n6970), 
	.B1(\fifo_from_fft/fifo_cell9/data_out/N35 ), 
	.B0(\fifo_from_fft/fifo_cell8/data_out/N35 ), 
	.A1(n4530), 
	.A0(n4536));
   XOR2X1TS U5683 (.Y(n6971), 
	.B(n6970), 
	.A(n6969));
   XOR2X1TS U5684 (.Y(n6972), 
	.B(n6971), 
	.A(n6968));
   AOI22X1TS U5685 (.Y(n6973), 
	.B1(\fifo_from_fft/fifo_cell13/data_out/N35 ), 
	.B0(\fifo_from_fft/fifo_cell1/data_out/N35 ), 
	.A1(n4578), 
	.A0(n4506));
   AOI22X1TS U5686 (.Y(n6974), 
	.B1(\fifo_from_fft/fifo_cell6/data_out/N35 ), 
	.B0(\fifo_from_fft/fifo_cell5/data_out/N35 ), 
	.A1(n4548), 
	.A0(n4554));
   XOR2X1TS U5687 (.Y(n6975), 
	.B(n6974), 
	.A(n6973));
   AOI22X1TS U5688 (.Y(n6976), 
	.B1(\fifo_from_fft/fifo_cell4/data_out/N35 ), 
	.B0(\fifo_from_fft/fifo_cell3/data_out/N35 ), 
	.A1(n4560), 
	.A0(n4566));
   XOR2X1TS U5689 (.Y(n6977), 
	.B(n6976), 
	.A(n4572));
   XOR2X1TS U5690 (.Y(n6978), 
	.B(n6977), 
	.A(n6975));
   AOI22X1TS U5691 (.Y(n6979), 
	.B1(\fifo_from_fft/fifo_cell15/data_out/N35 ), 
	.B0(\fifo_from_fft/fifo_cell10/data_out/N35 ), 
	.A1(n4524), 
	.A0(n4494));
   XOR2X1TS U5692 (.Y(n6980), 
	.B(n6979), 
	.A(n6978));
   XOR2X1TS U5693 (.Y(n6981), 
	.B(n6980), 
	.A(n6972));
   OAI21X1TS U5694 (.Y(n4580), 
	.B0(FE_OFN724_n4643), 
	.A1(n6981), 
	.A0(\fifo_from_fft/fifo_cell15/reg_gtok/token ));
   NOR3X1TS U5695 (.Y(n6982), 
	.C(\fifo_from_fir/fifo_cell0/controller/write_enable ), 
	.B(n7217), 
	.A(\fifo_from_fir/fifo_cell0/controller/valid_read ));
   AOI31X1TS U5696 (.Y(\fifo_from_fir/fifo_cell0/reg_ptok/N29 ), 
	.B0(\fifo_from_fir/hold[0] ), 
	.A2(n6982), 
	.A1(n3776), 
	.A0(\fifo_from_fir/fifo_cell0/data_out/N35 ));
   NOR3BX1TS U5697 (.Y(n3952), 
	.C(n3851), 
	.B(n8805), 
	.AN(\fifo_to_fft/hang[0] ));
   NOR3BX1TS U5698 (.Y(n4127), 
	.C(n4026), 
	.B(n8784), 
	.AN(\fifo_to_fir/hang[0] ));
   NOR2BX1TS U5699 (.Y(\add_x_22_2/carry[30] ), 
	.B(n7253), 
	.AN(\add_x_22_2/carry[29] ));
   XNOR2X1TS U5700 (.Y(\router/addr_calc/fir_read_calc/counter/N75 ), 
	.B(\add_x_22_2/carry[29] ), 
	.A(n7253));
   NOR3X1TS U5701 (.Y(n6983), 
	.C(\fifo_from_fft/fifo_cell8/controller/write_enable ), 
	.B(n7490), 
	.A(\fifo_from_fft/fifo_cell8/controller/valid_read ));
   AOI31X1TS U5702 (.Y(n4474), 
	.B0(\fifo_from_fft/hold[8] ), 
	.A2(n6983), 
	.A1(\fifo_from_fft/fifo_cell8/data_out/N35 ), 
	.A0(FE_OFN233_n4531));
   NOR3X1TS U5703 (.Y(n6984), 
	.C(\fifo_to_fir/fifo_cell5/controller/write_enable ), 
	.B(n7420), 
	.A(\fifo_to_fir/fifo_cell5/controller/valid_read ));
   AOI31X1TS U5704 (.Y(n4036), 
	.B0(\fifo_to_fir/hold[5] ), 
	.A2(n6984), 
	.A1(\fifo_to_fir/fifo_cell5/data_out/N35 ), 
	.A0(n7424));
   NOR3X1TS U5705 (.Y(n6985), 
	.C(\fifo_to_fft/fifo_cell11/controller/write_enable ), 
	.B(n7271), 
	.A(\fifo_to_fft/fifo_cell11/controller/valid_read ));
   AOI31X1TS U5706 (.Y(n3873), 
	.B0(\fifo_to_fft/hold[11] ), 
	.A2(n6985), 
	.A1(\fifo_to_fft/fifo_cell11/data_out/N35 ), 
	.A0(n3907));
   NOR3X1TS U5707 (.Y(n6986), 
	.C(\fifo_to_fir/fifo_cell12/controller/write_enable ), 
	.B(n7370), 
	.A(\fifo_to_fir/fifo_cell12/controller/valid_read ));
   AOI31X1TS U5708 (.Y(n4050), 
	.B0(\fifo_to_fir/hold[12] ), 
	.A2(n6986), 
	.A1(\fifo_to_fir/fifo_cell12/data_out/N35 ), 
	.A0(n7374));
   NOR3X1TS U5709 (.Y(n6987), 
	.C(\fifo_to_fft/fifo_cell13/controller/write_enable ), 
	.B(n7252), 
	.A(\fifo_to_fft/fifo_cell13/controller/valid_read ));
   AOI31X1TS U5710 (.Y(n3877), 
	.B0(\fifo_to_fft/hold[13] ), 
	.A2(n6987), 
	.A1(n7255), 
	.A0(\fifo_to_fft/fifo_cell13/data_out/N35 ));
   NOR3X1TS U5711 (.Y(n6988), 
	.C(\fifo_to_fir/fifo_cell14/controller/write_enable ), 
	.B(n7356), 
	.A(\fifo_to_fir/fifo_cell14/controller/valid_read ));
   AOI31X1TS U5712 (.Y(n4054), 
	.B0(\fifo_to_fir/hold[14] ), 
	.A2(n6988), 
	.A1(n4067), 
	.A0(\fifo_to_fir/fifo_cell14/data_out/N35 ));
   NOR2X1TS U5713 (.Y(n6989), 
	.B(n3764), 
	.A(n3763));
   OAI2BB2XLTS U5714 (.Y(n6990), 
	.B1(FE_OFN799_n7619), 
	.B0(FE_OFN682_n8050), 
	.A1N(n6989), 
	.A0N(n3767));
   OAI211X1TS U5715 (.Y(n5383), 
	.C0(n6990), 
	.B0(n9463), 
	.A1(n3760), 
	.A0(FE_OFN682_n8050));
   XOR2X1TS U5716 (.Y(n6991), 
	.B(n7199), 
	.A(\add_x_22_5/carry[31] ));
   AOI22X1TS U5717 (.Y(n6992), 
	.B1(n7198), 
	.B0(FE_OFN940_n3486), 
	.A1(n6991), 
	.A0(FE_OFN939_n3487));
   NAND2X1TS U5718 (.Y(\router/addr_calc/iir_write_calc/counter/N209 ), 
	.B(n6992), 
	.A(FE_OFN1295_iir_enable));
   AOI222XLTS U5719 (.Y(n3752), 
	.C1(fir_data_in[1]), 
	.C0(FE_OFN749_n3722), 
	.B1(FE_MDBN4_), 
	.B0(FE_OFN759_n3721), 
	.A1(\router/data_cntl/data_in[1] ), 
	.A0(FE_OFN770_n3720));
   AOI222XLTS U5720 (.Y(n3730), 
	.C1(fir_data_in[23]), 
	.C0(FE_OFN751_n3722), 
	.B1(fft_data_in[23]), 
	.B0(FE_OFN761_n3721), 
	.A1(\router/data_cntl/data_in[23] ), 
	.A0(FE_OFN772_n3720));
   AOI222XLTS U5721 (.Y(n3719), 
	.C1(FE_MDBN2_), 
	.C0(FE_OFN745_n3722), 
	.B1(FE_MDBN14_), 
	.B0(n3721), 
	.A1(\router/data_cntl/data_in[31] ), 
	.A0(FE_OFN766_n3720));
   AOI31X1TS U5722 (.Y(n6993), 
	.B0(n3715), 
	.A2(\router/fir_read_done ), 
	.A1(n9406), 
	.A0(FE_OFN976_n9462));
   NOR4X2TS U5723 (.Y(n4829), 
	.D(n6993), 
	.C(n7603), 
	.B(from_fir_empty), 
	.A(FE_OFN839_n7619));
   AOI22X1TS U5724 (.Y(n6994), 
	.B1(\fifo_from_fir/fifo_cell4/data_out/N35 ), 
	.B0(\fifo_from_fir/fifo_cell3/data_out/N35 ), 
	.A1(n4746), 
	.A0(n4752));
   AOI22X1TS U5725 (.Y(n6995), 
	.B1(\fifo_from_fir/fifo_cell6/data_out/N35 ), 
	.B0(\fifo_from_fir/fifo_cell5/data_out/N35 ), 
	.A1(n4734), 
	.A0(n4740));
   AOI22X1TS U5726 (.Y(n6996), 
	.B1(\fifo_from_fir/fifo_cell13/data_out/N35 ), 
	.B0(\fifo_from_fir/fifo_cell1/data_out/N35 ), 
	.A1(n4764), 
	.A0(n4692));
   XOR2X1TS U5727 (.Y(n6997), 
	.B(n6995), 
	.A(n6996));
   XOR2X1TS U5728 (.Y(n6998), 
	.B(n6994), 
	.A(n4758));
   XOR2X1TS U5729 (.Y(n6999), 
	.B(n6998), 
	.A(n6997));
   AOI22X1TS U5730 (.Y(n7000), 
	.B1(\fifo_from_fir/fifo_cell15/data_out/N35 ), 
	.B0(\fifo_from_fir/fifo_cell10/data_out/N35 ), 
	.A1(n4710), 
	.A0(n4680));
   AOI22X1TS U5731 (.Y(n7001), 
	.B1(\fifo_from_fir/fifo_cell12/data_out/N35 ), 
	.B0(\fifo_from_fir/fifo_cell11/data_out/N35 ), 
	.A1(n4698), 
	.A0(n4704));
   AOI22X1TS U5732 (.Y(n7002), 
	.B1(\fifo_from_fir/fifo_cell9/data_out/N35 ), 
	.B0(\fifo_from_fir/fifo_cell8/data_out/N35 ), 
	.A1(n4716), 
	.A0(n4722));
   AOI22X1TS U5733 (.Y(n7003), 
	.B1(\fifo_from_fir/fifo_cell14/data_out/N35 ), 
	.B0(\fifo_from_fir/fifo_cell7/data_out/N35 ), 
	.A1(n4728), 
	.A0(n4686));
   XOR2X1TS U5734 (.Y(n7004), 
	.B(n7002), 
	.A(n7001));
   XOR2X1TS U5735 (.Y(n7005), 
	.B(n7004), 
	.A(n7003));
   XOR2X1TS U5736 (.Y(n7006), 
	.B(n7000), 
	.A(n6999));
   XOR2X1TS U5737 (.Y(n7007), 
	.B(n7006), 
	.A(n7005));
   OAI21X1TS U5738 (.Y(n4766), 
	.B0(FE_OFN742_n4829), 
	.A1(n7007), 
	.A0(\fifo_from_fir/fifo_cell15/reg_gtok/token ));
   AND4X1TS U5739 (.Y(n7008), 
	.D(instruction[28]), 
	.C(instruction[0]), 
	.B(instruction[29]), 
	.A(instruction[27]));
   NAND4BX1TS U5740 (.Y(n7009), 
	.D(acc_bypass), 
	.C(n7008), 
	.B(instruction[26]), 
	.AN(n3458));
   AOI211X1TS U5741 (.Y(\router/pla_top/N60 ), 
	.C0(n7009), 
	.B0(n3456), 
	.A1(instruction[2]), 
	.A0(n3455));
   OAI21X1TS U5742 (.Y(n7010), 
	.B0(to_fft_empty), 
	.A1(n3476), 
	.A0(n3477));
   AND3X1TS U5743 (.Y(\router/data_cntl/N133 ), 
	.C(n7010), 
	.B(n9434), 
	.A(FE_OFN1217_n3478));
   NOR3X1TS U5744 (.Y(n7011), 
	.C(\fifo_from_fft/fifo_cell0/controller/write_enable ), 
	.B(n7222), 
	.A(\fifo_from_fft/fifo_cell0/controller/valid_read ));
   AOI31X1TS U5745 (.Y(\fifo_from_fft/fifo_cell0/reg_ptok/N29 ), 
	.B0(\fifo_from_fft/hold[0] ), 
	.A2(n7011), 
	.A1(n3796), 
	.A0(\fifo_from_fft/fifo_cell0/data_out/N35 ));
   NOR3X1TS U5746 (.Y(n7012), 
	.C(\fifo_to_fir/fifo_cell0/controller/write_enable ), 
	.B(n7227), 
	.A(\fifo_to_fir/fifo_cell0/controller/valid_read ));
   AOI31X1TS U5747 (.Y(\fifo_to_fir/fifo_cell0/reg_ptok/N29 ), 
	.B0(\fifo_to_fir/hold[0] ), 
	.A2(n7012), 
	.A1(n4136), 
	.A0(\fifo_to_fir/fifo_cell0/data_out/N35 ));
   NOR3X1TS U5748 (.Y(n7013), 
	.C(\fifo_to_fft/fifo_cell0/controller/write_enable ), 
	.B(n7232), 
	.A(\fifo_to_fft/fifo_cell0/controller/valid_read ));
   AOI31X1TS U5749 (.Y(\fifo_to_fft/fifo_cell0/reg_ptok/N29 ), 
	.B0(\fifo_to_fft/hold[0] ), 
	.A2(n7013), 
	.A1(n3961), 
	.A0(\fifo_to_fft/fifo_cell0/data_out/N35 ));
   CLKINVX2TS U5774 (.Y(n7014), 
	.A(\router/addr_calc/iir_write_calc/counter/hold ));
   INVX2TS U5775 (.Y(n7015), 
	.A(\router/addr_calc/N63 ));
   INVX2TS U5776 (.Y(n7016), 
	.A(\router/addr_calc/N95 ));
   INVX1TS U5777 (.Y(n7017), 
	.A(\router/addr_calc/N9 ));
   INVX2TS U5778 (.Y(n7018), 
	.A(\router/addr_calc/N99 ));
   INVX2TS U5779 (.Y(n7019), 
	.A(\router/addr_calc/fft_write_calc/counter/hold ));
   INVXLTS U5780 (.Y(n7020), 
	.A(\router/addr_calc/fir_write_calc/counter/hold ));
   INVXLTS U5781 (.Y(n7021), 
	.A(\router/addr_calc/fft_read_calc/counter/hold ));
   INVX2TS U5782 (.Y(n7022), 
	.A(\router/addr_calc/fir_read_calc/counter/hold ));
   INVX2TS U5783 (.Y(n7023), 
	.A(\router/addr_calc/fir_read_calc/counter/hold ));
   NAND4X1TS U5787 (.Y(n521), 
	.D(n3707), 
	.C(n3840), 
	.B(n2633), 
	.A(n2634));
   NOR2BX1TS U5795 (.Y(n7056), 
	.B(n9384), 
	.AN(n8027));
   NOR2BX1TS U5796 (.Y(n7057), 
	.B(n9384), 
	.AN(n8037));
   NOR2BX1TS U5797 (.Y(n7058), 
	.B(n9384), 
	.AN(n8026));
   NOR2BX1TS U5798 (.Y(n7059), 
	.B(n9384), 
	.AN(n8036));
   NOR2BX1TS U5799 (.Y(n7060), 
	.B(n9385), 
	.AN(n8025));
   NOR2BX1TS U5800 (.Y(n7061), 
	.B(n9385), 
	.AN(n8035));
   NOR2BX1TS U5801 (.Y(n7062), 
	.B(n9385), 
	.AN(n8024));
   NOR2BX1TS U5802 (.Y(n7063), 
	.B(n9385), 
	.AN(n8011));
   NOR2BX1TS U5803 (.Y(n7064), 
	.B(n9381), 
	.AN(n8018));
   NOR2BX1TS U5804 (.Y(n7065), 
	.B(n9381), 
	.AN(n8015));
   NOR2BX1TS U5805 (.Y(n7066), 
	.B(n9381), 
	.AN(n8042));
   NOR2BX1TS U5806 (.Y(n7067), 
	.B(n9382), 
	.AN(n8041));
   NOR2BX1TS U5807 (.Y(n7068), 
	.B(n9382), 
	.AN(n8017));
   NOR2BX1TS U5808 (.Y(n7069), 
	.B(n9382), 
	.AN(n8013));
   NOR2BX1TS U5809 (.Y(n7070), 
	.B(n9382), 
	.AN(n8040));
   NOR2BX1TS U5810 (.Y(n7071), 
	.B(n9383), 
	.AN(n8029));
   NOR2BX1TS U5811 (.Y(n7072), 
	.B(n9383), 
	.AN(n8039));
   NOR2BX1TS U5812 (.Y(n7073), 
	.B(n9383), 
	.AN(n8028));
   NOR2BX1TS U5813 (.Y(n7074), 
	.B(n9383), 
	.AN(n8038));
   NOR2BX1TS U5814 (.Y(n7075), 
	.B(n9381), 
	.AN(n8014));
   NOR2BX1TS U5815 (.Y(n7076), 
	.B(n9386), 
	.AN(n8034));
   NOR2BX1TS U5816 (.Y(n7077), 
	.B(n9386), 
	.AN(n8023));
   NOR2BX1TS U5817 (.Y(n7078), 
	.B(n9386), 
	.AN(n8033));
   NOR2BX1TS U5818 (.Y(n7079), 
	.B(n9386), 
	.AN(n8022));
   NOR2BX1TS U5819 (.Y(n7080), 
	.B(n9388), 
	.AN(n8030));
   NOR2BX1TS U5820 (.Y(n7081), 
	.B(n9388), 
	.AN(n8019));
   NOR2BX1TS U5821 (.Y(n7082), 
	.B(n9388), 
	.AN(n8016));
   NOR2BX1TS U5822 (.Y(n7083), 
	.B(n9388), 
	.AN(n8012));
   NOR2BX1TS U5823 (.Y(n7084), 
	.B(n9387), 
	.AN(n8032));
   NOR2BX1TS U5824 (.Y(n7085), 
	.B(n9387), 
	.AN(n8021));
   NOR2BX1TS U5825 (.Y(n7086), 
	.B(n9387), 
	.AN(n8031));
   NOR2BX1TS U5826 (.Y(n7087), 
	.B(n9387), 
	.AN(n8020));
   INVX1TS U5827 (.Y(n8715), 
	.A(FE_OFN174_n8054));
   INVX1TS U5828 (.Y(n8716), 
	.A(FE_OFN174_n8054));
   CLKINVX2TS U5829 (.Y(n8713), 
	.A(FE_OFN173_n8054));
   INVX1TS U5830 (.Y(n8717), 
	.A(FE_OFN174_n8054));
   INVX1TS U5831 (.Y(n8718), 
	.A(n8054));
   CLKINVX2TS U5832 (.Y(n8714), 
	.A(FE_OFN174_n8054));
   CLKINVX2TS U5833 (.Y(n8712), 
	.A(FE_OFN173_n8054));
   INVX1TS U5834 (.Y(n8378), 
	.A(FE_OFN509_n8055));
   INVX1TS U5835 (.Y(n8379), 
	.A(FE_OFN510_n8055));
   INVX1TS U5836 (.Y(n8382), 
	.A(FE_OFN510_n8055));
   INVX1TS U5837 (.Y(n8384), 
	.A(FE_OFN508_n8055));
   INVX1TS U5838 (.Y(n8381), 
	.A(FE_OFN510_n8055));
   INVX1TS U5839 (.Y(n8383), 
	.A(FE_OFN508_n8055));
   INVX1TS U5840 (.Y(n8380), 
	.A(FE_OFN510_n8055));
   INVXLTS U5841 (.Y(n8719), 
	.A(FE_OFN173_n8054));
   INVX1TS U5842 (.Y(n8377), 
	.A(FE_OFN509_n8055));
   INVX1TS U5843 (.Y(n7366), 
	.A(n4072));
   INVX1TS U5844 (.Y(n7256), 
	.A(n3897));
   INVX2TS U5845 (.Y(n7255), 
	.A(n3897));
   INVX2TS U5846 (.Y(n7365), 
	.A(n4072));
   INVX2TS U5847 (.Y(n7374), 
	.A(n4077));
   INVX2TS U5848 (.Y(n7265), 
	.A(n3902));
   CLKINVX1TS U5849 (.Y(n7286), 
	.A(n3917));
   CLKINVX1TS U5850 (.Y(n7395), 
	.A(n4092));
   INVX2TS U5851 (.Y(n7394), 
	.A(n4092));
   INVX2TS U5852 (.Y(n7285), 
	.A(n3917));
   INVX2TS U5853 (.Y(n7295), 
	.A(n3922));
   INVX2TS U5854 (.Y(n7404), 
	.A(n4097));
   INVX2TS U5855 (.Y(n7315), 
	.A(n3937));
   INVX2TS U5856 (.Y(n7424), 
	.A(n4112));
   CLKINVX1TS U5857 (.Y(n7316), 
	.A(n3937));
   CLKINVX1TS U5858 (.Y(n7425), 
	.A(n4112));
   INVX1TS U5859 (.Y(n8143), 
	.A(FE_OFN665_n8053));
   INVX1TS U5860 (.Y(n8144), 
	.A(n8053));
   INVX1TS U5861 (.Y(n8141), 
	.A(FE_OFN665_n8053));
   CLKINVX2TS U5862 (.Y(n8140), 
	.A(FE_OFN665_n8053));
   INVX1TS U5863 (.Y(n8142), 
	.A(FE_OFN665_n8053));
   CLKINVX2TS U5864 (.Y(n8139), 
	.A(FE_OFN664_n8053));
   INVX1TS U5865 (.Y(n8473), 
	.A(FE_OFN326_n8056));
   INVX1TS U5866 (.Y(n8474), 
	.A(FE_OFN326_n8056));
   INVX1TS U5867 (.Y(n8480), 
	.A(FE_OFN326_n8056));
   INVX1TS U5868 (.Y(n8479), 
	.A(FE_OFN326_n8056));
   INVX1TS U5869 (.Y(n8475), 
	.A(FE_OFN325_n8056));
   INVX1TS U5870 (.Y(n8478), 
	.A(FE_OFN325_n8056));
   INVX1TS U5871 (.Y(n8476), 
	.A(FE_OFN325_n8056));
   CLKINVX2TS U5872 (.Y(n8138), 
	.A(FE_OFN664_n8053));
   INVX1TS U5873 (.Y(n8477), 
	.A(n8056));
   CLKINVX1TS U5874 (.Y(n8145), 
	.A(n8053));
   INVX1TS U5875 (.Y(n8790), 
	.A(n8057));
   CLKINVX2TS U5876 (.Y(n8789), 
	.A(FE_OFN734_n8057));
   INVX1TS U5877 (.Y(n8787), 
	.A(FE_OFN733_n8057));
   CLKINVX1TS U5878 (.Y(n8876), 
	.A(FE_OFN679_n8050));
   CLKINVX1TS U5879 (.Y(n8843), 
	.A(n8052));
   INVX1TS U5880 (.Y(n8811), 
	.A(FE_OFN731_n8058));
   INVX2TS U5881 (.Y(n7444), 
	.A(n4128));
   INVX1TS U5882 (.Y(n8808), 
	.A(FE_OFN729_n8058));
   CLKINVX1TS U5883 (.Y(n8842), 
	.A(FE_OFN697_n8052));
   INVX2TS U5884 (.Y(n7335), 
	.A(n3953));
   CLKINVX2TS U5885 (.Y(n8810), 
	.A(FE_OFN730_n8058));
   CLKINVX1TS U5886 (.Y(n8875), 
	.A(FE_OFN679_n8050));
   CLKINVX1TS U5887 (.Y(n7445), 
	.A(n4128));
   CLKINVX2TS U5888 (.Y(n7236), 
	.A(n3883));
   INVX1TS U5889 (.Y(n7616), 
	.A(n4057));
   INVX1TS U5890 (.Y(n7615), 
	.A(n4057));
   INVX1TS U5891 (.Y(n7614), 
	.A(n4057));
   INVXLTS U5892 (.Y(n8845), 
	.A(FE_OFN698_n8052));
   AND4X1TS U5893 (.Y(n8057), 
	.D(n7608), 
	.C(n9465), 
	.B(\router/fir_put_req_reg ), 
	.A(n3715));
   CLKINVX1TS U5894 (.Y(n8873), 
	.A(FE_OFN680_n8050));
   INVXLTS U5895 (.Y(n8878), 
	.A(FE_OFN682_n8050));
   INVX1TS U5896 (.Y(n7617), 
	.A(n4057));
   CLKINVX1TS U5897 (.Y(n7336), 
	.A(n3953));
   CLKINVX1TS U5898 (.Y(n8840), 
	.A(FE_OFN696_n8052));
   CLKINVX2TS U5899 (.Y(n7345), 
	.A(n4058));
   INVX2TS U5900 (.Y(n7608), 
	.A(n3474));
   INVX1TS U5901 (.Y(n8870), 
	.A(n8050));
   INVX1TS U5902 (.Y(n8837), 
	.A(n8052));
   CLKINVX1TS U5903 (.Y(n8841), 
	.A(FE_OFN697_n8052));
   CLKINVX1TS U5904 (.Y(n8874), 
	.A(FE_OFN680_n8050));
   CLKINVX1TS U5905 (.Y(n9378), 
	.A(FE_OFN718_n8051));
   OR2X2TS U5906 (.Y(n4057), 
	.B(FE_OFN687_n4134), 
	.A(FE_OFN800_n7619));
   CLKINVX2TS U5907 (.Y(n9372), 
	.A(FE_OFN717_n8051));
   CLKINVX2TS U5908 (.Y(n9376), 
	.A(FE_OFN718_n8051));
   CLKINVX2TS U5909 (.Y(n9370), 
	.A(n8051));
   CLKINVX2TS U5910 (.Y(n9377), 
	.A(FE_OFN718_n8051));
   CLKINVX2TS U5911 (.Y(n9371), 
	.A(n8051));
   CLKINVX2TS U5912 (.Y(n9373), 
	.A(FE_OFN717_n8051));
   CLKINVX1TS U5913 (.Y(n9375), 
	.A(FE_OFN718_n8051));
   CLKINVX1TS U5914 (.Y(n9374), 
	.A(FE_OFN717_n8051));
   INVX1TS U5915 (.Y(n7971), 
	.A(n7967));
   INVX1TS U5916 (.Y(n7970), 
	.A(n7967));
   CLKAND2X2TS U5917 (.Y(n5580), 
	.B(\mips/mips/accfullinstruction[25] ), 
	.A(FE_OFN711_n4207));
   INVX1TS U5918 (.Y(n7968), 
	.A(n7967));
   CLKAND2X2TS U5919 (.Y(n5581), 
	.B(\mips/mips/accfullinstruction[24] ), 
	.A(FE_OFN710_n4207));
   CLKAND2X2TS U5920 (.Y(n5582), 
	.B(\mips/mips/accfullinstruction[23] ), 
	.A(FE_OFN713_n4207));
   CLKAND2X2TS U5921 (.Y(n5583), 
	.B(\mips/mips/accfullinstruction[22] ), 
	.A(FE_OFN711_n4207));
   INVX1TS U5922 (.Y(n7969), 
	.A(n7967));
   OR2X2TS U5923 (.Y(n8051), 
	.B(\mips/mips/a/N49 ), 
	.A(\mips/mips/a/countflag ));
   INVX1TS U5924 (.Y(n7965), 
	.A(n7962));
   INVX1TS U5925 (.Y(n7964), 
	.A(n7962));
   INVX1TS U5926 (.Y(n7963), 
	.A(n7962));
   INVX1TS U5927 (.Y(n7966), 
	.A(n7962));
   INVX2TS U5928 (.Y(n7593), 
	.A(n4756));
   CLKINVX2TS U5929 (.Y(n7490), 
	.A(n4534));
   INVX2TS U5930 (.Y(n7369), 
	.A(n4076));
   INVX2TS U5931 (.Y(n7568), 
	.A(n4726));
   INVX2TS U5932 (.Y(n7280), 
	.A(n3916));
   CLKINVX2TS U5933 (.Y(n7514), 
	.A(n4564));
   CLKINVX2TS U5934 (.Y(n7232), 
	.A(n3820));
   CLKINVX1TS U5935 (.Y(n7470), 
	.A(n4510));
   INVX2TS U5936 (.Y(n7414), 
	.A(n4106));
   INVX2TS U5937 (.Y(n7464), 
	.A(n4504));
   CLKAND2X2TS U5938 (.Y(n5600), 
	.B(\mips/mips/accfullinstruction[5] ), 
	.A(FE_OFN711_n4207));
   INVX2TS U5939 (.Y(n7409), 
	.A(n4101));
   INVX2TS U5940 (.Y(n7563), 
	.A(n4720));
   INVX2TS U5941 (.Y(n7270), 
	.A(n3906));
   INVX2TS U5942 (.Y(n7493), 
	.A(n4540));
   INVX2TS U5943 (.Y(n7484), 
	.A(n4528));
   CLKINVX1TS U5944 (.Y(n7356), 
	.A(n4066));
   INVX2TS U5945 (.Y(n7553), 
	.A(n4708));
   INVX2TS U5946 (.Y(n7275), 
	.A(n3911));
   INVX2TS U5947 (.Y(n7558), 
	.A(n4714));
   INVX2TS U5948 (.Y(n7379), 
	.A(n4081));
   INVX2TS U5949 (.Y(n7459), 
	.A(n4498));
   CLKINVX1TS U5950 (.Y(n7480), 
	.A(n4522));
   INVX2TS U5951 (.Y(n7548), 
	.A(n4702));
   INVX2TS U5952 (.Y(n7260), 
	.A(n3901));
   INVX2TS U5953 (.Y(n7399), 
	.A(n4096));
   CLKINVX1TS U5954 (.Y(n7361), 
	.A(n4071));
   INVX2TS U5955 (.Y(n7384), 
	.A(n4086));
   CLKINVX2TS U5956 (.Y(n7370), 
	.A(n4076));
   CLKINVX1TS U5957 (.Y(n7242), 
	.A(n3886));
   INVX2TS U5958 (.Y(n7251), 
	.A(n3896));
   INVX1TS U5959 (.Y(n7252), 
	.A(n3896));
   CLKINVX1TS U5960 (.Y(n7594), 
	.A(n4756));
   INVX2TS U5961 (.Y(n7469), 
	.A(n4510));
   CLKINVX2TS U5962 (.Y(n7380), 
	.A(n4081));
   INVX2TS U5963 (.Y(n7573), 
	.A(n4732));
   CLKAND2X2TS U5964 (.Y(n5579), 
	.B(\mips/mips/accfullinstruction[26] ), 
	.A(n7977));
   CLKINVX1TS U5965 (.Y(n7321), 
	.A(n3941));
   CLKINVX2TS U5966 (.Y(n7261), 
	.A(n3901));
   INVX2TS U5967 (.Y(n7598), 
	.A(n4762));
   INVX2TS U5968 (.Y(n7216), 
	.A(n3774));
   CLKINVX2TS U5969 (.Y(n7385), 
	.A(n4086));
   INVX1TS U5970 (.Y(n7311), 
	.A(n3936));
   INVX2TS U5971 (.Y(n7246), 
	.A(n3891));
   CLKINVX1TS U5972 (.Y(n7430), 
	.A(n4116));
   INVX2TS U5973 (.Y(n7538), 
	.A(n4690));
   INVX2TS U5974 (.Y(n7474), 
	.A(n4516));
   CLKINVX2TS U5975 (.Y(n7271), 
	.A(n3906));
   INVX2TS U5976 (.Y(n7533), 
	.A(n4684));
   INVX2TS U5977 (.Y(n7241), 
	.A(n3886));
   CLKINVX2TS U5978 (.Y(n7390), 
	.A(n4091));
   CLKAND2X2TS U5979 (.Y(n5577), 
	.B(\mips/mips/accfullinstruction[28] ), 
	.A(n7977));
   INVX2TS U5980 (.Y(n7301), 
	.A(n3926));
   INVX1TS U5981 (.Y(n7485), 
	.A(n4528));
   INVX1TS U5982 (.Y(n7420), 
	.A(n4111));
   INVX2TS U5983 (.Y(n7543), 
	.A(n4696));
   INVX2TS U5984 (.Y(n7489), 
	.A(n4534));
   INVX2TS U5985 (.Y(n7389), 
	.A(n4091));
   CLKINVX2TS U5986 (.Y(n7291), 
	.A(n3921));
   INVX2TS U5987 (.Y(n7276), 
	.A(n3911));
   CLKINVX2TS U5988 (.Y(n7400), 
	.A(n4096));
   CLKINVX2TS U5989 (.Y(n7415), 
	.A(n4106));
   INVX2TS U5990 (.Y(n7281), 
	.A(n3916));
   CLKINVX2TS U5991 (.Y(n7410), 
	.A(n4101));
   CLKAND2X2TS U5992 (.Y(n5578), 
	.B(\mips/mips/accfullinstruction[27] ), 
	.A(n7977));
   INVX2TS U5993 (.Y(n7330), 
	.A(n3951));
   INVX2TS U5994 (.Y(n7226), 
	.A(n3809));
   INVX2TS U5995 (.Y(n7325), 
	.A(n3946));
   INVX2TS U5996 (.Y(n7449), 
	.A(n4131));
   INVX2TS U5997 (.Y(n7429), 
	.A(n4116));
   INVX2TS U5998 (.Y(n7340), 
	.A(n3956));
   CLKINVX2TS U5999 (.Y(n7574), 
	.A(n4732));
   INVX2TS U6000 (.Y(n7498), 
	.A(n4546));
   INVX2TS U6001 (.Y(n7231), 
	.A(n3820));
   CLKINVX2TS U6002 (.Y(n7569), 
	.A(n4726));
   INVX2TS U6003 (.Y(n7588), 
	.A(n4750));
   INVX2TS U6004 (.Y(n7320), 
	.A(n3941));
   INVX2TS U6005 (.Y(n7503), 
	.A(n4552));
   CLKINVX1TS U6006 (.Y(n7475), 
	.A(n4516));
   CLKINVX1TS U6007 (.Y(n7554), 
	.A(n4708));
   INVX2TS U6008 (.Y(n7310), 
	.A(n3936));
   INVX2TS U6009 (.Y(n7583), 
	.A(n4744));
   CLKINVX2TS U6010 (.Y(n7564), 
	.A(n4720));
   INVX2TS U6011 (.Y(n7439), 
	.A(n4126));
   INVX2TS U6012 (.Y(n7454), 
	.A(n4492));
   CLKINVX2TS U6013 (.Y(n7579), 
	.A(n4738));
   CLKINVX2TS U6014 (.Y(n7227), 
	.A(n3809));
   INVX2TS U6015 (.Y(n7528), 
	.A(n4678));
   CLKINVX2TS U6016 (.Y(n7509), 
	.A(n4558));
   CLKINVX1TS U6017 (.Y(n7247), 
	.A(n3891));
   CLKINVX1TS U6018 (.Y(n7559), 
	.A(n4714));
   INVX2TS U6019 (.Y(n7513), 
	.A(n4564));
   CLKINVX1TS U6020 (.Y(n7544), 
	.A(n4696));
   CLKINVX2TS U6021 (.Y(n7504), 
	.A(n4552));
   INVX2TS U6022 (.Y(n7434), 
	.A(n4121));
   INVX2TS U6023 (.Y(n7419), 
	.A(n4111));
   INVX2TS U6024 (.Y(n7508), 
	.A(n4558));
   INVX2TS U6025 (.Y(n7355), 
	.A(n4066));
   INVX2TS U6026 (.Y(n7479), 
	.A(n4522));
   CLKINVX2TS U6027 (.Y(n7584), 
	.A(n4744));
   INVX2TS U6028 (.Y(n7578), 
	.A(n4738));
   CLKINVX1TS U6029 (.Y(n7549), 
	.A(n4702));
   CLKINVX2TS U6030 (.Y(n7499), 
	.A(n4546));
   INVX2TS U6031 (.Y(n7290), 
	.A(n3921));
   INVX1TS U6032 (.Y(n7589), 
	.A(n4750));
   INVX2TS U6033 (.Y(n7300), 
	.A(n3926));
   CLKINVX2TS U6034 (.Y(n7360), 
	.A(n4071));
   CLKINVX2TS U6035 (.Y(n7494), 
	.A(n4540));
   INVX2TS U6036 (.Y(n7203), 
	.A(FE_OFN973_n7207));
   INVX1TS U6037 (.Y(n7977), 
	.A(n3456));
   CLKINVX2TS U6038 (.Y(n7306), 
	.A(n3931));
   CLKINVX1TS U6039 (.Y(n7351), 
	.A(n4061));
   INVX2TS U6040 (.Y(n7305), 
	.A(n3931));
   AND2XLTS U6041 (.Y(n5576), 
	.B(\mips/mips/accfullinstruction[29] ), 
	.A(n4205));
   AND2XLTS U6042 (.Y(n5574), 
	.B(\mips/mips/accfullinstruction[31] ), 
	.A(n4205));
   AND2XLTS U6043 (.Y(n5575), 
	.B(\mips/mips/accfullinstruction[30] ), 
	.A(n4205));
   INVX2TS U6044 (.Y(n7518), 
	.A(n4570));
   CLKINVX1TS U6045 (.Y(n7524), 
	.A(n4576));
   INVX2TS U6046 (.Y(n7221), 
	.A(n3794));
   CLKINVX2TS U6047 (.Y(n9463), 
	.A(FE_OFN793_n7619));
   CLKINVX2TS U6048 (.Y(n9545), 
	.A(FE_OFN807_n7619));
   CLKINVX2TS U6049 (.Y(n9464), 
	.A(FE_OFN789_n7619));
   CLKINVX2TS U6050 (.Y(n9546), 
	.A(FE_OFN785_n7619));
   CLKINVX2TS U6051 (.Y(n9543), 
	.A(FE_OFN815_n7619));
   INVX1TS U6052 (.Y(n7519), 
	.A(n4570));
   CLKINVX2TS U6053 (.Y(n9544), 
	.A(FE_OFN812_n7619));
   INVX2TS U6054 (.Y(n7350), 
	.A(n4061));
   INVX2TS U6055 (.Y(n7523), 
	.A(n4576));
   CLKINVX2TS U6056 (.Y(n9525), 
	.A(FE_OFN811_n7619));
   CLKINVX2TS U6057 (.Y(n9521), 
	.A(FE_OFN832_n7619));
   CLKINVX2TS U6058 (.Y(n9509), 
	.A(FE_OFN795_n7619));
   CLKINVX2TS U6059 (.Y(n9528), 
	.A(FE_OFN821_n7619));
   CLKINVX2TS U6060 (.Y(n9508), 
	.A(FE_OFN796_n7619));
   CLKINVX2TS U6061 (.Y(n9488), 
	.A(FE_OFN799_n7619));
   CLKINVX2TS U6062 (.Y(n9516), 
	.A(FE_OFN790_n7619));
   CLKINVX2TS U6063 (.Y(n9520), 
	.A(FE_OFN791_n7619));
   CLKINVX2TS U6064 (.Y(n9522), 
	.A(FE_OFN824_n7619));
   CLKINVX2TS U6065 (.Y(n9524), 
	.A(FE_OFN787_n7619));
   CLKINVX2TS U6066 (.Y(n9517), 
	.A(FE_OFN826_n7619));
   CLKINVX2TS U6067 (.Y(n9547), 
	.A(FE_OFN784_n7619));
   CLKINVX2TS U6068 (.Y(n9531), 
	.A(FE_OFN778_n7619));
   CLKINVX2TS U6069 (.Y(n9493), 
	.A(FE_OFN811_n7619));
   CLKINVX2TS U6070 (.Y(n9512), 
	.A(FE_OFN815_n7619));
   CLKINVX2TS U6071 (.Y(n9530), 
	.A(FE_OFN822_n7619));
   CLKINVX2TS U6072 (.Y(n9510), 
	.A(FE_OFN795_n7619));
   CLKINVX2TS U6073 (.Y(n9529), 
	.A(FE_OFN808_n7619));
   CLKINVX2TS U6074 (.Y(n9526), 
	.A(FE_OFN816_n7619));
   CLKINVX2TS U6075 (.Y(n9515), 
	.A(FE_OFN784_n7619));
   CLKINVX2TS U6076 (.Y(n9511), 
	.A(FE_OFN793_n7619));
   CLKINVX2TS U6077 (.Y(n9518), 
	.A(FE_OFN842_n7619));
   CLKINVX2TS U6078 (.Y(n9479), 
	.A(FE_OFN813_n7619));
   CLKINVX2TS U6079 (.Y(n9478), 
	.A(FE_OFN797_n7619));
   CLKINVX2TS U6080 (.Y(n9495), 
	.A(FE_OFN810_n7619));
   CLKINVX2TS U6081 (.Y(n9474), 
	.A(FE_OFN790_n7619));
   CLKINVX2TS U6082 (.Y(n9519), 
	.A(FE_OFN792_n7619));
   CLKINVX2TS U6083 (.Y(n9491), 
	.A(FE_OFN801_n7619));
   CLKINVX2TS U6084 (.Y(n9523), 
	.A(FE_OFN802_n7619));
   CLKINVX2TS U6085 (.Y(n9492), 
	.A(FE_OFN777_n7619));
   CLKINVX2TS U6086 (.Y(n9477), 
	.A(FE_OFN797_n7619));
   CLKINVX2TS U6087 (.Y(n9527), 
	.A(FE_OFN814_n7619));
   CLKINVX2TS U6088 (.Y(n9489), 
	.A(FE_OFN786_n7619));
   CLKINVX2TS U6089 (.Y(n7606), 
	.A(n8059));
   INVX2TS U6090 (.Y(n7207), 
	.A(n3472));
   CLKINVX2TS U6091 (.Y(n9501), 
	.A(FE_OFN798_n7619));
   CLKINVX2TS U6092 (.Y(n9539), 
	.A(FE_OFN781_n7619));
   CLKINVX2TS U6093 (.Y(n9502), 
	.A(FE_OFN814_n7619));
   CLKINVX2TS U6094 (.Y(n9540), 
	.A(FE_OFN818_n7619));
   CLKINVX2TS U6095 (.Y(n9541), 
	.A(FE_OFN830_n7619));
   CLKINVX2TS U6096 (.Y(n9535), 
	.A(FE_OFN800_n7619));
   CLKINVX2TS U6097 (.Y(n9467), 
	.A(FE_OFN831_n7619));
   CLKINVX2TS U6098 (.Y(n9500), 
	.A(FE_OFN805_n7619));
   CLKINVX2TS U6099 (.Y(n9466), 
	.A(FE_OFN833_n7619));
   CLKINVX2TS U6100 (.Y(n9507), 
	.A(FE_OFN830_n7619));
   CLKINVX2TS U6101 (.Y(n9542), 
	.A(FE_OFN783_n7619));
   CLKINVX2TS U6102 (.Y(n9503), 
	.A(FE_OFN823_n7619));
   CLKINVX2TS U6103 (.Y(n9471), 
	.A(FE_OFN827_n7619));
   CLKINVX2TS U6104 (.Y(n9468), 
	.A(FE_OFN815_n7619));
   CLKINVX2TS U6105 (.Y(n9532), 
	.A(FE_OFN834_n7619));
   CLKINVX2TS U6106 (.Y(n9533), 
	.A(FE_OFN826_n7619));
   CLKINVX2TS U6107 (.Y(n9534), 
	.A(FE_OFN819_n7619));
   CLKINVX2TS U6108 (.Y(n9506), 
	.A(FE_OFN780_n7619));
   CLKINVX2TS U6109 (.Y(n9505), 
	.A(FE_OFN793_n7619));
   CLKINVX2TS U6110 (.Y(n9504), 
	.A(FE_OFN777_n7619));
   CLKINVX2TS U6111 (.Y(n9496), 
	.A(FE_OFN834_n7619));
   CLKINVX2TS U6112 (.Y(n9498), 
	.A(FE_OFN801_n7619));
   CLKINVX2TS U6113 (.Y(n9499), 
	.A(FE_OFN838_n7619));
   CLKINVX1TS U6114 (.Y(n9434), 
	.A(FE_OFN974_n9462));
   CLKINVX2TS U6115 (.Y(n9415), 
	.A(FE_OFN993_n9431));
   CLKINVX2TS U6116 (.Y(n9442), 
	.A(FE_OFN982_n9462));
   CLKINVX4TS U6117 (.Y(fft_enable), 
	.A(FE_OFN983_n9462));
   CLKINVX2TS U6118 (.Y(n9414), 
	.A(FE_OFN987_n9431));
   NAND3XLTS U6119 (.Y(n8059), 
	.C(FE_OFN1286_iir_enable), 
	.B(FE_OFN991_n9431), 
	.A(FE_OFN979_n9462));
   INVX2TS U6120 (.Y(n7610), 
	.A(FE_OFN1285_router_ram_read_enable_reg));
   CLKINVX1TS U6121 (.Y(n9443), 
	.A(FE_OFN982_n9462));
   CLKINVX1TS U6122 (.Y(n9439), 
	.A(FE_OFN975_n9462));
   INVX1TS U6123 (.Y(n9445), 
	.A(FE_OFN983_n9462));
   CLKINVX2TS U6124 (.Y(n7611), 
	.A(FE_OFN1285_router_ram_read_enable_reg));
   CLKINVX1TS U6125 (.Y(n9440), 
	.A(FE_OFN975_n9462));
   INVX1TS U6126 (.Y(n9444), 
	.A(FE_OFN983_n9462));
   INVXLTS U6127 (.Y(n9391), 
	.A(iir_enable));
   CLKINVX2TS U6128 (.Y(n9447), 
	.A(FE_OFN984_n9462));
   CLKINVX2TS U6129 (.Y(n9420), 
	.A(FE_OFN992_n9431));
   CLKINVX1TS U6130 (.Y(n9417), 
	.A(FE_OFN993_n9431));
   CLKINVX1TS U6131 (.Y(n9416), 
	.A(FE_OFN992_n9431));
   INVX2TS U6132 (.Y(n7603), 
	.A(\router/fir_get_req_reg ));
   CLKINVX2TS U6133 (.Y(n9421), 
	.A(FE_OFN992_n9431));
   INVX2TS U6134 (.Y(n7211), 
	.A(\router/fir_read_done ));
   CLKINVX2TS U6135 (.Y(n9446), 
	.A(FE_OFN984_n9462));
   CLKINVX2TS U6136 (.Y(n9470), 
	.A(FE_OFN812_n7619));
   CLKINVX1TS U6137 (.Y(n7960), 
	.A(n4458));
   INVX1TS U6138 (.Y(n7527), 
	.A(n7525));
   CLKINVX1TS U6139 (.Y(n7157), 
	.A(n7155));
   CLKINVX1TS U6140 (.Y(n7151), 
	.A(n7149));
   CLKINVX1TS U6141 (.Y(n7162), 
	.A(n7161));
   INVX1TS U6142 (.Y(n7403), 
	.A(n7401));
   INVX1TS U6144 (.Y(n7393), 
	.A(n7391));
   CLKINVX2TS U6145 (.Y(n7398), 
	.A(n7396));
   CLKINVX1TS U6146 (.Y(n7378), 
	.A(n7376));
   CLKINVX1TS U6147 (.Y(n7502), 
	.A(n7500));
   INVX1TS U6148 (.Y(n7166), 
	.A(n7164));
   INVX1TS U6149 (.Y(n7154), 
	.A(n7152));
   CLKINVX2TS U6150 (.Y(n7160), 
	.A(n7158));
   CLKINVX1TS U6151 (.Y(n7130), 
	.A(n7128));
   CLKINVX1TS U6152 (.Y(n7373), 
	.A(n7371));
   CLKINVX1TS U6153 (.Y(n7497), 
	.A(n7495));
   CLKINVX1TS U6154 (.Y(n7168), 
	.A(n7167));
   CLKINVX1TS U6155 (.Y(n7147), 
	.A(n7146));
   CLKINVX1TS U6156 (.Y(n7387), 
	.A(n7386));
   CLKINVX1TS U6157 (.Y(n7511), 
	.A(n7510));
   CLKINVX2TS U6158 (.Y(n7192), 
	.A(n7191));
   CLKINVX1TS U6159 (.Y(n7174), 
	.A(n7173));
   INVX1TS U6160 (.Y(n7186), 
	.A(n7185));
   CLKINVX1TS U6161 (.Y(n7141), 
	.A(n7140));
   CLKINVX1TS U6162 (.Y(n7382), 
	.A(n7381));
   CLKINVX1TS U6163 (.Y(n7506), 
	.A(n7505));
   CLKINVX1TS U6165 (.Y(n7199), 
	.A(n7197));
   CLKINVX1TS U6166 (.Y(n7136), 
	.A(n7134));
   CLKINVX1TS U6167 (.Y(n7442), 
	.A(n7441));
   CLKINVX1TS U6168 (.Y(n7189), 
	.A(n7188));
   CLKINVX1TS U6169 (.Y(n7224), 
	.A(n7223));
   CLKINVX2TS U6170 (.Y(n7522), 
	.A(n7520));
   CLKINVX1TS U6171 (.Y(n7089), 
	.A(n7088));
   CLKINVX1TS U6172 (.Y(n7422), 
	.A(n7421));
   CLKINVX1TS U6173 (.Y(n7546), 
	.A(n7545));
   CLKINVX1TS U6174 (.Y(n7132), 
	.A(n7131));
   CLKINVX1TS U6175 (.Y(n7183), 
	.A(n7182));
   CLKINVX1TS U6176 (.Y(n7541), 
	.A(n7540));
   CLKINVX1TS U6177 (.Y(n7096), 
	.A(n7094));
   CLKINVX1TS U6178 (.Y(n7591), 
	.A(n7590));
   CLKINVX1TS U6179 (.Y(n7417), 
	.A(n7416));
   CLKINVX1TS U6180 (.Y(n7472), 
	.A(n7471));
   CLKINVX1TS U6181 (.Y(n7138), 
	.A(n7137));
   CLKINVX1TS U6182 (.Y(n7234), 
	.A(n7233));
   CLKINVX1TS U6183 (.Y(n7177), 
	.A(n7176));
   CLKINVX1TS U6184 (.Y(n7101), 
	.A(n7100));
   CLKINVX1TS U6185 (.Y(n7596), 
	.A(n7595));
   CLKINVX1TS U6186 (.Y(n7412), 
	.A(n7411));
   CLKINVX1TS U6187 (.Y(n7477), 
	.A(n7476));
   CLKINVX1TS U6188 (.Y(n7536), 
	.A(n7535));
   CLKINVX1TS U6189 (.Y(n7145), 
	.A(n7143));
   CLKINVX1TS U6190 (.Y(n7566), 
	.A(n7565));
   INVX1TS U6191 (.Y(n7289), 
	.A(n7287));
   CLKINVX1TS U6192 (.Y(n7109), 
	.A(n7108));
   CLKINVX1TS U6193 (.Y(n7309), 
	.A(n7307));
   CLKINVX1TS U6194 (.Y(n7209), 
	.A(n7208));
   CLKINVX1TS U6195 (.Y(n7304), 
	.A(n7302));
   CLKINVX1TS U6196 (.Y(n7205), 
	.A(n7204));
   CLKINVX1TS U6197 (.Y(n7104), 
	.A(n7103));
   INVX2TS U6198 (.Y(n7258), 
	.A(n7257));
   CLKINVX2TS U6199 (.Y(n7263), 
	.A(n7262));
   CLKINVX1TS U6200 (.Y(n7437), 
	.A(n7436));
   CLKINVX1TS U6201 (.Y(n7561), 
	.A(n7560));
   CLKINVX1TS U6202 (.Y(n7329), 
	.A(n7327));
   CLKINVX1TS U6203 (.Y(n7115), 
	.A(n7114));
   CLKINVX1TS U6204 (.Y(n7571), 
	.A(n7570));
   CLKINVX1TS U6205 (.Y(n7201), 
	.A(n7200));
   CLKINVX1TS U6206 (.Y(n7447), 
	.A(n7446));
   CLKINVX1TS U6207 (.Y(n7318), 
	.A(n7317));
   CLKINVX1TS U6208 (.Y(n7359), 
	.A(n7357));
   INVX1TS U6209 (.Y(n7517), 
	.A(n7515));
   CLKINVX1TS U6210 (.Y(n7432), 
	.A(n7431));
   CLKINVX1TS U6211 (.Y(n7214), 
	.A(n7213));
   CLKINVX1TS U6212 (.Y(n7354), 
	.A(n7352));
   CLKINVX1TS U6213 (.Y(n7556), 
	.A(n7555));
   CLKINVX1TS U6214 (.Y(n7098), 
	.A(n7097));
   INVX1TS U6215 (.Y(n7279), 
	.A(n7277));
   CLKINVX2TS U6216 (.Y(n7284), 
	.A(n7282));
   CLKINVX1TS U6217 (.Y(n7334), 
	.A(n7332));
   CLKINVX1TS U6218 (.Y(n7576), 
	.A(n7575));
   CLKINVX1TS U6219 (.Y(n7121), 
	.A(n7120));
   CLKINVX1TS U6220 (.Y(n7324), 
	.A(n7322));
   CLKINVX1TS U6221 (.Y(n7299), 
	.A(n7297));
   CLKINVX1TS U6222 (.Y(n7452), 
	.A(n7451));
   CLKINVX1TS U6223 (.Y(n7338), 
	.A(n7337));
   CLKINVX1TS U6224 (.Y(n7195), 
	.A(n7194));
   CLKINVX1TS U6225 (.Y(n7219), 
	.A(n7218));
   CLKINVX1TS U6226 (.Y(n7313), 
	.A(n7312));
   CLKINVX1TS U6227 (.Y(n7427), 
	.A(n7426));
   CLKINVX1TS U6228 (.Y(n7092), 
	.A(n7091));
   INVX1TS U6229 (.Y(n7269), 
	.A(n7267));
   CLKINVX1TS U6230 (.Y(n7581), 
	.A(n7580));
   CLKINVX1TS U6231 (.Y(n7551), 
	.A(n7550));
   INVX1TS U6232 (.Y(n7274), 
	.A(n7272));
   CLKINVX1TS U6233 (.Y(n7457), 
	.A(n7456));
   CLKINVX1TS U6234 (.Y(n7126), 
	.A(n7125));
   CLKINVX1TS U6235 (.Y(n7343), 
	.A(n7342));
   CLKINVX1TS U6236 (.Y(n7408), 
	.A(n7406));
   CLKINVX1TS U6237 (.Y(n7239), 
	.A(n7238));
   CLKINVX1TS U6238 (.Y(n7172), 
	.A(n7170));
   CLKINVX1TS U6239 (.Y(n7113), 
	.A(n7111));
   CLKINVX1TS U6240 (.Y(n7532), 
	.A(n7530));
   CLKINVX1TS U6241 (.Y(n7294), 
	.A(n7292));
   INVX1TS U6242 (.Y(n7180), 
	.A(n7179));
   INVX2TS U6243 (.Y(n1161), 
	.A(\fifo_from_fft/fifo_cell9/data_out/N9 ));
   INVX2TS U6244 (.Y(n2569), 
	.A(\fifo_from_fir/fifo_cell15/data_out/N9 ));
   INVX2TS U6245 (.Y(n1289), 
	.A(\fifo_from_fft/fifo_cell11/data_out/N9 ));
   INVX2TS U6246 (.Y(n1353), 
	.A(\fifo_from_fft/fifo_cell12/data_out/N9 ));
   INVX2TS U6247 (.Y(n2441), 
	.A(\fifo_from_fir/fifo_cell13/data_out/N9 ));
   INVX2TS U6248 (.Y(n1417), 
	.A(\fifo_from_fft/fifo_cell13/data_out/N9 ));
   INVX2TS U6249 (.Y(n2377), 
	.A(\fifo_from_fir/fifo_cell12/data_out/N9 ));
   INVX2TS U6250 (.Y(n1225), 
	.A(\fifo_from_fft/fifo_cell10/data_out/N9 ));
   INVX2TS U6251 (.Y(n1097), 
	.A(\fifo_from_fft/fifo_cell8/data_out/N9 ));
   INVX2TS U6252 (.Y(n2505), 
	.A(\fifo_from_fir/fifo_cell14/data_out/N9 ));
   INVX2TS U6253 (.Y(n2313), 
	.A(\fifo_from_fir/fifo_cell11/data_out/N9 ));
   INVX1TS U6254 (.Y(n585), 
	.A(\fifo_from_fft/fifo_cell0/data_out/N9 ));
   INVX2TS U6255 (.Y(n1481), 
	.A(\fifo_from_fft/fifo_cell14/data_out/N9 ));
   INVX2TS U6256 (.Y(n1673), 
	.A(\fifo_from_fir/fifo_cell1/data_out/N9 ));
   INVX2TS U6257 (.Y(n1033), 
	.A(\fifo_from_fft/fifo_cell7/data_out/N9 ));
   INVX2TS U6258 (.Y(n2249), 
	.A(\fifo_from_fir/fifo_cell10/data_out/N9 ));
   INVX2TS U6259 (.Y(n649), 
	.A(\fifo_from_fft/fifo_cell1/data_out/N9 ));
   INVX1TS U6260 (.Y(n1609), 
	.A(\fifo_from_fir/fifo_cell0/data_out/N9 ));
   INVX2TS U6261 (.Y(n1737), 
	.A(\fifo_from_fir/fifo_cell2/data_out/N9 ));
   INVX2TS U6262 (.Y(n1545), 
	.A(\fifo_from_fft/fifo_cell15/data_out/N9 ));
   INVX2TS U6263 (.Y(n969), 
	.A(\fifo_from_fft/fifo_cell6/data_out/N9 ));
   INVX2TS U6264 (.Y(n2185), 
	.A(\fifo_from_fir/fifo_cell9/data_out/N9 ));
   INVX2TS U6265 (.Y(n713), 
	.A(\fifo_from_fft/fifo_cell2/data_out/N9 ));
   INVX2TS U6266 (.Y(n1801), 
	.A(\fifo_from_fir/fifo_cell3/data_out/N9 ));
   INVX2TS U6267 (.Y(n905), 
	.A(\fifo_from_fft/fifo_cell5/data_out/N9 ));
   INVX2TS U6268 (.Y(n1865), 
	.A(\fifo_from_fir/fifo_cell4/data_out/N9 ));
   INVX2TS U6269 (.Y(n2121), 
	.A(\fifo_from_fir/fifo_cell8/data_out/N9 ));
   INVX2TS U6270 (.Y(n1929), 
	.A(\fifo_from_fir/fifo_cell5/data_out/N9 ));
   INVX2TS U6271 (.Y(n841), 
	.A(\fifo_from_fft/fifo_cell4/data_out/N9 ));
   INVX2TS U6272 (.Y(n2057), 
	.A(\fifo_from_fir/fifo_cell7/data_out/N9 ));
   INVX2TS U6273 (.Y(n777), 
	.A(\fifo_from_fft/fifo_cell3/data_out/N9 ));
   INVX2TS U6275 (.Y(n1993), 
	.A(\fifo_from_fir/fifo_cell6/data_out/N9 ));
   INVX2TS U6277 (.Y(n137), 
	.A(\router/addr_calc/N191 ));
   INVX2TS U6278 (.Y(n9431), 
	.A(n9615));
   INVX2TS U6279 (.Y(n9462), 
	.A(n9614));
   INVXLTS U6538 (.Y(n7119), 
	.A(n7117));
   INVXLTS U6539 (.Y(n7212), 
	.A(\router/fir_read_done ));
   INVXLTS U6540 (.Y(n7217), 
	.A(n3774));
   INVXLTS U6541 (.Y(n7222), 
	.A(n3794));
   INVXLTS U6542 (.Y(n7230), 
	.A(n7228));
   INVXLTS U6543 (.Y(n7237), 
	.A(n3883));
   INVXLTS U6544 (.Y(n7245), 
	.A(n7243));
   CLKINVX2TS U6545 (.Y(n7250), 
	.A(n7248));
   INVXLTS U6546 (.Y(n7266), 
	.A(n3902));
   INVXLTS U6548 (.Y(n7326), 
	.A(n3946));
   INVXLTS U6549 (.Y(n7331), 
	.A(n3951));
   INVXLTS U6550 (.Y(n7341), 
	.A(n3956));
   INVXLTS U6551 (.Y(n7346), 
	.A(n4058));
   CLKINVX2TS U6552 (.Y(n7349), 
	.A(n7347));
   CLKINVX2TS U6553 (.Y(n7364), 
	.A(n7362));
   INVXLTS U6554 (.Y(n7375), 
	.A(n4077));
   INVXLTS U6555 (.Y(n7405), 
	.A(n4097));
   INVXLTS U6556 (.Y(n7435), 
	.A(n4121));
   INVXLTS U6557 (.Y(n7440), 
	.A(n4126));
   INVXLTS U6558 (.Y(n7450), 
	.A(n4131));
   INVXLTS U6559 (.Y(n7455), 
	.A(n4492));
   INVXLTS U6560 (.Y(n7460), 
	.A(n4498));
   INVXLTS U6561 (.Y(n7463), 
	.A(n7461));
   INVXLTS U6562 (.Y(n7465), 
	.A(n4504));
   INVXLTS U6563 (.Y(n7468), 
	.A(n7466));
   CLKINVX2TS U6564 (.Y(n7483), 
	.A(n7481));
   INVXLTS U6565 (.Y(n7488), 
	.A(n7486));
   INVXLTS U6566 (.Y(n7529), 
	.A(n4678));
   INVXLTS U6567 (.Y(n7534), 
	.A(n4684));
   INVXLTS U6568 (.Y(n7539), 
	.A(n4690));
   INVXLTS U6569 (.Y(n7587), 
	.A(n7585));
   INVXLTS U6570 (.Y(n7599), 
	.A(n4762));
   INVXLTS U6571 (.Y(n7602), 
	.A(n7600));
   INVXLTS U6572 (.Y(n7607), 
	.A(n8059));
   INVXLTS U6573 (.Y(n7609), 
	.A(n3474));
   INVX2TS U6574 (.Y(n7618), 
	.A(FE_OFN1447_reset));
   INVX2TS U6575 (.Y(n7619), 
	.A(n7618));
   AND3X2TS U6576 (.Y(n8050), 
	.C(n3465), 
	.B(n9514), 
	.A(FE_OFN1451_acc_fir_put));
   AND3X2TS U6577 (.Y(n8052), 
	.C(n3477), 
	.B(n9513), 
	.A(FE_OFN1449_acc_fft_put));
   INVX2TS U6651 (.Y(n7953), 
	.A(n4025));
   OR2X2TS U6653 (.Y(n7962), 
	.B(FE_OFN741_n4829), 
	.A(FE_OFN828_n7619));
   OR2X2TS U6654 (.Y(n7967), 
	.B(FE_OFN728_n4643), 
	.A(FE_OFN847_n7619));
   INVX2TS U6655 (.Y(n7973), 
	.A(n7972));
   INVX2TS U6656 (.Y(n7976), 
	.A(n7972));
   INVX2TS U6657 (.Y(n7975), 
	.A(n7972));
   INVX2TS U6658 (.Y(n7974), 
	.A(n7972));
   XOR2X1TS U6659 (.Y(\router/addr_calc/fft_read_calc/counter/N77 ), 
	.B(n7488), 
	.A(\add_x_22_0/carry[31] ));
   XOR2X1TS U6661 (.Y(\router/addr_calc/fft_write_calc/counter/N77 ), 
	.B(\router/addr_calc/fft_write_calc/count[31] ), 
	.A(\add_x_22_1/carry[31] ));
   XOR2X1TS U6663 (.Y(\router/addr_calc/fir_read_calc/counter/N77 ), 
	.B(n7250), 
	.A(\add_x_22_2/carry[31] ));
   XOR2X1TS U6665 (.Y(\router/addr_calc/fir_write_calc/counter/N77 ), 
	.B(n7119), 
	.A(\add_x_22_3/carry[31] ));
   INVX2TS U6684 (.Y(n8872), 
	.A(FE_OFN680_n8050));
   INVX2TS U6689 (.Y(n8839), 
	.A(FE_OFN697_n8052));
   INVX2TS U6741 (.Y(n9537), 
	.A(FE_OFN785_n7619));
   INVX2TS U6742 (.Y(n9536), 
	.A(FE_OFN779_n7619));
   INVX2TS U6743 (.Y(n9538), 
	.A(FE_OFN781_n7619));
   INVX2TS U6744 (.Y(n9390), 
	.A(iir_enable));
   INVX2TS U6745 (.Y(n9389), 
	.A(FE_OFN1286_iir_enable));
   INVX2TS U6766 (.Y(fir_enable), 
	.A(FE_OFN986_n9431));
   INVX2TS U6777 (.Y(n9475), 
	.A(FE_OFN816_n7619));
   INVX2TS U6778 (.Y(n8809), 
	.A(FE_OFN731_n8058));
   INVX2TS U6779 (.Y(n8788), 
	.A(FE_OFN734_n8057));
   INVX2TS U6782 (.Y(n9476), 
	.A(FE_OFN819_n7619));
   INVX2TS U6785 (.Y(n8791), 
	.A(FE_OFN732_n8057));
   INVX2TS U6786 (.Y(n8812), 
	.A(FE_OFN730_n8058));
   INVX2TS U6790 (.Y(n9472), 
	.A(FE_OFN789_n7619));
   INVX2TS U6791 (.Y(n9469), 
	.A(FE_OFN799_n7619));
   INVX2TS U6792 (.Y(n9473), 
	.A(FE_OFN777_n7619));
   AND2X2TS U6793 (.Y(n5603), 
	.B(\mips/mips/accfullinstruction[2] ), 
	.A(n4207));
   AND2X2TS U6794 (.Y(n5602), 
	.B(\mips/mips/accfullinstruction[3] ), 
	.A(FE_OFN709_n4207));
   INVX2TS U6811 (.Y(n9448), 
	.A(FE_OFN984_n9462));
   INVX2TS U6812 (.Y(n9413), 
	.A(FE_OFN989_n9431));
   INVX2TS U6813 (.Y(n9449), 
	.A(FE_OFN984_n9462));
   INVX2TS U6822 (.Y(n9490), 
	.A(FE_OFN842_n7619));
   INVX2TS U6823 (.Y(n9494), 
	.A(FE_OFN823_n7619));
   INVX2TS U6841 (.Y(n9484), 
	.A(FE_OFN809_n7619));
   INVX2TS U6842 (.Y(n9483), 
	.A(FE_OFN806_n7619));
   INVX2TS U6843 (.Y(n9482), 
	.A(FE_OFN824_n7619));
   INVX2TS U6844 (.Y(n9481), 
	.A(FE_OFN825_n7619));
   OAI22XLTS U6845 (.Y(n6233), 
	.B1(n3755), 
	.B0(n3841), 
	.A1(n3843), 
	.A0(n3754));
   INVX2TS U6847 (.Y(n9438), 
	.A(FE_OFN975_n9462));
   INVX2TS U6848 (.Y(n9419), 
	.A(FE_OFN993_n9431));
   INVX2TS U6851 (.Y(n9437), 
	.A(FE_OFN980_n9462));
   INVX2TS U6852 (.Y(n9436), 
	.A(FE_OFN980_n9462));
   INVX2TS U6855 (.Y(n9418), 
	.A(FE_OFN993_n9431));
   INVX2TS U6856 (.Y(n9441), 
	.A(FE_OFN975_n9462));
   INVX2TS U6871 (.Y(n9487), 
	.A(FE_OFN788_n7619));
   INVX2TS U6872 (.Y(n9486), 
	.A(FE_OFN817_n7619));
endmodule

