library verilog;
use verilog.vl_types.all;
entity CLKINVX4TS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end CLKINVX4TS;
