library verilog;
use verilog.vl_types.all;
entity TIELOTS is
    port(
        Y               : out    vl_logic
    );
end TIELOTS;
