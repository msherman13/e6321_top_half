library verilog;
use verilog.vl_types.all;
entity udp_mux is
    // This module cannot be connected to from
    // VHDL because it has unnamed ports.
end udp_mux;
