library verilog;
use verilog.vl_types.all;
entity DLY1X1TS is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end DLY1X1TS;
